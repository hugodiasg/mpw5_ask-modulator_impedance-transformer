magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< pwell >>
rect -191 1002 191 1088
rect -191 -1002 -105 1002
rect 105 -1002 191 1002
rect -191 -1088 191 -1002
<< psubdiff >>
rect -165 1028 -51 1062
rect -17 1028 17 1062
rect 51 1028 165 1062
rect -165 935 -131 1028
rect 131 935 165 1028
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect -165 -1028 -131 -935
rect 131 -1028 165 -935
rect -165 -1062 -51 -1028
rect -17 -1062 17 -1028
rect 51 -1062 165 -1028
<< psubdiffcont >>
rect -51 1028 -17 1062
rect 17 1028 51 1062
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect -51 -1062 -17 -1028
rect 17 -1062 51 -1028
<< xpolycontact >>
rect -35 500 35 932
rect -35 -932 35 -500
<< xpolyres >>
rect -35 -500 35 500
<< locali >>
rect -165 1028 -51 1062
rect -17 1028 17 1062
rect 51 1028 165 1062
rect -165 935 -131 1028
rect 131 1025 165 1028
rect 131 953 165 991
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect 131 881 165 901
rect 131 809 165 833
rect 131 737 165 765
rect 131 665 165 697
rect 131 595 165 629
rect 131 527 165 559
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect 131 459 165 487
rect 131 391 165 415
rect 131 323 165 343
rect 131 255 165 271
rect 131 187 165 199
rect 131 119 165 127
rect 131 51 165 55
rect 131 -55 165 -51
rect 131 -127 165 -119
rect 131 -199 165 -187
rect 131 -271 165 -255
rect 131 -343 165 -323
rect 131 -415 165 -391
rect 131 -487 165 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect 131 -559 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -665
rect 131 -765 165 -737
rect 131 -833 165 -809
rect 131 -901 165 -881
rect -165 -1028 -131 -935
rect 131 -991 165 -953
rect 131 -1028 165 -1025
rect -165 -1062 -51 -1028
rect -17 -1062 17 -1028
rect 51 -1062 165 -1028
<< viali >>
rect 131 991 165 1025
rect 131 935 165 953
rect -17 878 17 912
rect -17 806 17 840
rect -17 734 17 768
rect -17 662 17 696
rect -17 590 17 624
rect -17 518 17 552
rect 131 919 165 935
rect 131 867 165 881
rect 131 847 165 867
rect 131 799 165 809
rect 131 775 165 799
rect 131 731 165 737
rect 131 703 165 731
rect 131 663 165 665
rect 131 631 165 663
rect 131 561 165 593
rect 131 559 165 561
rect 131 493 165 521
rect 131 487 165 493
rect 131 425 165 449
rect 131 415 165 425
rect 131 357 165 377
rect 131 343 165 357
rect 131 289 165 305
rect 131 271 165 289
rect 131 221 165 233
rect 131 199 165 221
rect 131 153 165 161
rect 131 127 165 153
rect 131 85 165 89
rect 131 55 165 85
rect 131 -17 165 17
rect 131 -85 165 -55
rect 131 -89 165 -85
rect 131 -153 165 -127
rect 131 -161 165 -153
rect 131 -221 165 -199
rect 131 -233 165 -221
rect 131 -289 165 -271
rect 131 -305 165 -289
rect 131 -357 165 -343
rect 131 -377 165 -357
rect 131 -425 165 -415
rect 131 -449 165 -425
rect 131 -493 165 -487
rect -17 -553 17 -519
rect -17 -625 17 -591
rect -17 -697 17 -663
rect -17 -769 17 -735
rect -17 -841 17 -807
rect -17 -913 17 -879
rect 131 -521 165 -493
rect 131 -561 165 -559
rect 131 -593 165 -561
rect 131 -663 165 -631
rect 131 -665 165 -663
rect 131 -731 165 -703
rect 131 -737 165 -731
rect 131 -799 165 -775
rect 131 -809 165 -799
rect 131 -867 165 -847
rect 131 -881 165 -867
rect 131 -935 165 -919
rect 131 -953 165 -935
rect 131 -1025 165 -991
<< metal1 >>
rect 125 1025 171 1040
rect 125 991 131 1025
rect 165 991 171 1025
rect 125 953 171 991
rect -25 912 25 926
rect -25 878 -17 912
rect 17 878 25 912
rect -25 840 25 878
rect -25 806 -17 840
rect 17 806 25 840
rect -25 768 25 806
rect -25 734 -17 768
rect 17 734 25 768
rect -25 696 25 734
rect -25 662 -17 696
rect 17 662 25 696
rect -25 624 25 662
rect -25 590 -17 624
rect 17 590 25 624
rect -25 552 25 590
rect -25 518 -17 552
rect 17 518 25 552
rect -25 505 25 518
rect 125 919 131 953
rect 165 919 171 953
rect 125 881 171 919
rect 125 847 131 881
rect 165 847 171 881
rect 125 809 171 847
rect 125 775 131 809
rect 165 775 171 809
rect 125 737 171 775
rect 125 703 131 737
rect 165 703 171 737
rect 125 665 171 703
rect 125 631 131 665
rect 165 631 171 665
rect 125 593 171 631
rect 125 559 131 593
rect 165 559 171 593
rect 125 521 171 559
rect 125 487 131 521
rect 165 487 171 521
rect 125 449 171 487
rect 125 415 131 449
rect 165 415 171 449
rect 125 377 171 415
rect 125 343 131 377
rect 165 343 171 377
rect 125 305 171 343
rect 125 271 131 305
rect 165 271 171 305
rect 125 233 171 271
rect 125 199 131 233
rect 165 199 171 233
rect 125 161 171 199
rect 125 127 131 161
rect 165 127 171 161
rect 125 89 171 127
rect 125 55 131 89
rect 165 55 171 89
rect 125 17 171 55
rect 125 -17 131 17
rect 165 -17 171 17
rect 125 -55 171 -17
rect 125 -89 131 -55
rect 165 -89 171 -55
rect 125 -127 171 -89
rect 125 -161 131 -127
rect 165 -161 171 -127
rect 125 -199 171 -161
rect 125 -233 131 -199
rect 165 -233 171 -199
rect 125 -271 171 -233
rect 125 -305 131 -271
rect 165 -305 171 -271
rect 125 -343 171 -305
rect 125 -377 131 -343
rect 165 -377 171 -343
rect 125 -415 171 -377
rect 125 -449 131 -415
rect 165 -449 171 -415
rect 125 -487 171 -449
rect -25 -519 25 -505
rect -25 -553 -17 -519
rect 17 -553 25 -519
rect -25 -591 25 -553
rect -25 -625 -17 -591
rect 17 -625 25 -591
rect -25 -663 25 -625
rect -25 -697 -17 -663
rect 17 -697 25 -663
rect -25 -735 25 -697
rect -25 -769 -17 -735
rect 17 -769 25 -735
rect -25 -807 25 -769
rect -25 -841 -17 -807
rect 17 -841 25 -807
rect -25 -879 25 -841
rect -25 -913 -17 -879
rect 17 -913 25 -879
rect -25 -926 25 -913
rect 125 -521 131 -487
rect 165 -521 171 -487
rect 125 -559 171 -521
rect 125 -593 131 -559
rect 165 -593 171 -559
rect 125 -631 171 -593
rect 125 -665 131 -631
rect 165 -665 171 -631
rect 125 -703 171 -665
rect 125 -737 131 -703
rect 165 -737 171 -703
rect 125 -775 171 -737
rect 125 -809 131 -775
rect 165 -809 171 -775
rect 125 -847 171 -809
rect 125 -881 131 -847
rect 165 -881 171 -847
rect 125 -919 171 -881
rect 125 -953 131 -919
rect 165 -953 171 -919
rect 125 -991 171 -953
rect 125 -1025 131 -991
rect 165 -1025 171 -991
rect 125 -1040 171 -1025
<< properties >>
string FIXED_BBOX -148 -1045 148 1045
<< end >>
