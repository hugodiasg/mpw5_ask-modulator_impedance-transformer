magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< pwell >>
rect 6534 -7232 6994 -6980
<< mvpsubdiff >>
rect 6560 -7021 6968 -7006
rect 6560 -7191 6611 -7021
rect 6917 -7191 6968 -7021
rect 6560 -7206 6968 -7191
<< mvpsubdiffcont >>
rect 6611 -7191 6917 -7021
<< locali >>
rect 6568 -7017 6960 -7006
rect 6568 -7195 6603 -7017
rect 6925 -7195 6960 -7017
rect 6568 -7206 6960 -7195
<< viali >>
rect 6603 -7021 6925 -7017
rect 6603 -7191 6611 -7021
rect 6611 -7191 6917 -7021
rect 6917 -7191 6925 -7021
rect 6603 -7195 6925 -7191
<< metal1 >>
rect 6300 16598 9480 16640
rect 6300 16162 8868 16598
rect 9432 16162 9480 16598
rect 6300 16120 9480 16162
rect 7700 -1682 9360 -1640
rect 7700 -2758 7750 -1682
rect 8570 -2180 9360 -1682
rect 10360 -1662 11560 -1620
rect 10360 -2098 10968 -1662
rect 11532 -2098 11560 -1662
rect 10360 -2158 11560 -2098
rect 10360 -2160 10954 -2158
rect 8570 -2758 8680 -2180
rect 8860 -2580 10360 -2240
rect 7700 -2800 8680 -2758
rect 9960 -2800 10360 -2580
rect 6340 -4480 9760 -2800
rect 9880 -3360 10360 -2800
rect 9880 -3740 10660 -3360
rect 9880 -4480 10360 -3740
rect 9718 -4646 9884 -4572
rect 9720 -5160 9880 -4646
rect 6340 -5360 9880 -5160
rect 10480 -6765 10660 -3740
rect 6572 -7006 6956 -7000
rect 10480 -7006 10664 -6765
rect 6344 -7017 10664 -7006
rect 6344 -7195 6603 -7017
rect 6925 -7195 10664 -7017
rect 6344 -7206 10664 -7195
rect 6572 -7212 6956 -7206
<< via1 >>
rect 8868 16162 9432 16598
rect 7750 -2758 8570 -1682
rect 10968 -2098 11532 -1662
<< metal2 >>
rect 8820 16608 9480 16640
rect 8820 16152 8842 16608
rect 9458 16152 9480 16608
rect 8820 16120 9480 16152
rect 7700 -1640 8600 -1620
rect 7700 -1682 8660 -1640
rect 7700 -1712 7750 -1682
rect 8570 -1712 8660 -1682
rect 7700 -2728 7732 -1712
rect 8588 -2728 8660 -1712
rect 10920 -1662 11580 -1600
rect 10920 -2098 10968 -1662
rect 11532 -2098 11580 -1662
rect 10920 -2140 11580 -2098
rect 7700 -2758 7750 -2728
rect 8570 -2758 8660 -2728
rect 7700 -2820 8660 -2758
<< via2 >>
rect 8842 16598 9458 16608
rect 8842 16162 8868 16598
rect 8868 16162 9432 16598
rect 9432 16162 9458 16598
rect 8842 16152 9458 16162
rect 7732 -2728 7750 -1712
rect 7750 -2728 8570 -1712
rect 8570 -2728 8588 -1712
rect 10982 -2068 11518 -1692
<< metal3 >>
rect 8820 16612 9480 16640
rect 8820 16608 8878 16612
rect 9422 16608 9480 16612
rect 8820 16152 8842 16608
rect 9458 16152 9480 16608
rect 8820 16148 8878 16152
rect 9422 16148 9480 16152
rect 8820 16120 9480 16148
rect 7700 -1640 8600 -1620
rect 7700 -1708 8660 -1640
rect 7700 -2732 7728 -1708
rect 8592 -2732 8660 -1708
rect 10920 -1688 11580 -1600
rect 10920 -2072 10978 -1688
rect 11522 -2072 11580 -1688
rect 10920 -2140 11580 -2072
rect 7700 -2820 8660 -2732
<< via3 >>
rect 8878 16608 9422 16612
rect 8878 16152 9422 16608
rect 8878 16148 9422 16152
rect 7728 -1712 8592 -1708
rect 7728 -2728 7732 -1712
rect 7732 -2728 8588 -1712
rect 8588 -2728 8592 -1712
rect 7728 -2732 8592 -2728
rect 10978 -1692 11522 -1688
rect 10978 -2068 10982 -1692
rect 10982 -2068 11518 -1692
rect 11518 -2068 11522 -1692
rect 10978 -2072 11522 -2068
<< metal4 >>
rect 8820 16612 9480 16640
rect 8820 16498 8878 16612
rect 9422 16498 9480 16612
rect 8820 16262 8872 16498
rect 9428 16262 9480 16498
rect 8820 16148 8878 16262
rect 9422 16148 9480 16262
rect 8820 16120 9480 16148
rect 7020 9040 12260 9420
rect 7020 3840 12260 4260
rect 7700 -1640 8600 -329
rect 9220 -380 15380 1980
rect 7700 -1708 8660 -1640
rect 7700 -2732 7728 -1708
rect 8592 -2732 8660 -1708
rect 10920 -1688 11580 -1600
rect 10920 -1762 10978 -1688
rect 11522 -1762 11580 -1688
rect 10920 -1998 10972 -1762
rect 11528 -1998 11580 -1762
rect 10920 -2072 10978 -1998
rect 11522 -2072 11580 -1998
rect 10920 -2140 11580 -2072
rect 7700 -2820 8660 -2732
rect 13020 -6420 15380 -380
rect 13020 -8780 30458 -6420
<< via4 >>
rect 8872 16262 8878 16498
rect 8878 16262 9108 16498
rect 9192 16262 9422 16498
rect 9422 16262 9428 16498
rect 10972 -1998 10978 -1762
rect 10978 -1998 11208 -1762
rect 11292 -1998 11522 -1762
rect 11522 -1998 11528 -1762
<< metal5 >>
rect 8819 16644 11980 17562
rect 8816 16498 11980 16644
rect 8816 16262 8872 16498
rect 9108 16262 9192 16498
rect 9428 16262 11980 16498
rect 8816 16116 11980 16262
rect 8819 15200 11980 16116
rect 12640 17560 12940 17562
rect 13860 17560 15123 17562
rect 12640 15200 15123 17560
rect 8819 12219 11181 15200
rect 9200 12200 10400 12219
rect 10940 -1600 11580 -338
rect 10920 -1762 11580 -1600
rect 10920 -1998 10972 -1762
rect 11208 -1998 11292 -1762
rect 11528 -1998 11580 -1762
rect 10920 -2140 11580 -1998
<< rm5 >>
rect 11980 15200 12640 17562
use l0_0  l0_0_0
timestamp 1647143569
transform 1 0 -24400 0 1 -45638
box 39200 36838 63200 63200
use sky130_fd_pr__cap_mim_m3_2_97K3D8  sky130_fd_pr__cap_mim_m3_2_97K3D8_0
timestamp 1647143569
transform -1 0 9641 0 1 6632
box -2619 -7770 2641 7770
use sky130_fd_pr__nfet_g5v0d10v5_PWYS4E  sky130_fd_pr__nfet_g5v0d10v5_PWYS4E_0
timestamp 1647143569
transform 1 0 9796 0 1 -3646
box -268 -1118 268 1118
use sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN  sky130_fd_pr__res_xhigh_po_0p35_CTQ8XN_0
timestamp 1647143569
transform 0 1 9872 -1 0 -2093
box -191 -1088 191 1088
<< labels >>
flabel metal1 s 6344 -7206 6544 -7006 0 FreeSans 160 0 0 0 gnd
port 1 nsew
flabel metal1 s 6340 -5360 6540 -5160 0 FreeSans 160 0 0 0 in
port 2 nsew
flabel metal1 s 6340 -3040 6540 -2840 0 FreeSans 160 0 0 0 out
port 3 nsew
flabel metal1 s 6340 16440 6540 16640 0 FreeSans 160 0 0 0 vd
port 4 nsew
<< end >>
