magic
tech sky130A
timestamp 1647143569
<< metal4 >>
rect 26249 24899 27429 24950
rect 26249 23821 26300 24899
rect 27378 23821 27429 24899
rect 26249 18419 27429 23821
<< via4 >>
rect 26300 23821 27378 24899
<< metal5 >>
rect 19600 30419 31600 31600
rect 19600 29029 30209 30209
rect 19600 20780 20780 29029
rect 20990 27639 28819 28819
rect 20990 22170 22170 27639
rect 22380 26249 27429 27429
rect 22380 23560 23560 26249
rect 26249 24899 27429 26249
rect 26249 23821 26300 24899
rect 27378 23821 27429 24899
rect 26249 23770 27429 23821
rect 27639 23560 28819 27639
rect 22380 22380 28819 23560
rect 29029 22170 30209 29029
rect 20990 20990 30209 22170
rect 30419 20780 31600 30419
rect 19600 19600 31600 20780
<< end >>
