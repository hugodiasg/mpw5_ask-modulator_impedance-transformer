magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< metal4 >>
rect -2472 7084 2472 7279
rect -2472 6848 2216 7084
rect 2452 6848 2472 7084
rect -2472 6764 2472 6848
rect -2472 6528 2216 6764
rect 2452 6528 2472 6764
rect -2472 6444 2472 6528
rect -2472 6208 2216 6444
rect 2452 6208 2472 6444
rect -2472 6124 2472 6208
rect -2472 5888 2216 6124
rect 2452 5888 2472 6124
rect -2472 5804 2472 5888
rect -2472 5568 2216 5804
rect 2452 5568 2472 5804
rect -2472 5484 2472 5568
rect -2472 5248 2216 5484
rect 2452 5248 2472 5484
rect -2472 5164 2472 5248
rect -2472 4928 2216 5164
rect 2452 4928 2472 5164
rect -2472 4844 2472 4928
rect -2472 4608 2216 4844
rect 2452 4608 2472 4844
rect -2472 4524 2472 4608
rect -2472 4288 2216 4524
rect 2452 4288 2472 4524
rect -2472 4204 2472 4288
rect -2472 3968 2216 4204
rect 2452 3968 2472 4204
rect -2472 3884 2472 3968
rect -2472 3648 2216 3884
rect 2452 3648 2472 3884
rect -2472 3564 2472 3648
rect -2472 3328 2216 3564
rect 2452 3328 2472 3564
rect -2472 3244 2472 3328
rect -2472 3008 2216 3244
rect 2452 3008 2472 3244
rect -2472 2924 2472 3008
rect -2472 2688 2216 2924
rect 2452 2688 2472 2924
rect -2472 2493 2472 2688
rect -2472 2198 2472 2393
rect -2472 1962 2216 2198
rect 2452 1962 2472 2198
rect -2472 1878 2472 1962
rect -2472 1642 2216 1878
rect 2452 1642 2472 1878
rect -2472 1558 2472 1642
rect -2472 1322 2216 1558
rect 2452 1322 2472 1558
rect -2472 1238 2472 1322
rect -2472 1002 2216 1238
rect 2452 1002 2472 1238
rect -2472 918 2472 1002
rect -2472 682 2216 918
rect 2452 682 2472 918
rect -2472 598 2472 682
rect -2472 362 2216 598
rect 2452 362 2472 598
rect -2472 278 2472 362
rect -2472 42 2216 278
rect 2452 42 2472 278
rect -2472 -42 2472 42
rect -2472 -278 2216 -42
rect 2452 -278 2472 -42
rect -2472 -362 2472 -278
rect -2472 -598 2216 -362
rect 2452 -598 2472 -362
rect -2472 -682 2472 -598
rect -2472 -918 2216 -682
rect 2452 -918 2472 -682
rect -2472 -1002 2472 -918
rect -2472 -1238 2216 -1002
rect 2452 -1238 2472 -1002
rect -2472 -1322 2472 -1238
rect -2472 -1558 2216 -1322
rect 2452 -1558 2472 -1322
rect -2472 -1642 2472 -1558
rect -2472 -1878 2216 -1642
rect 2452 -1878 2472 -1642
rect -2472 -1962 2472 -1878
rect -2472 -2198 2216 -1962
rect 2452 -2198 2472 -1962
rect -2472 -2393 2472 -2198
rect -2472 -2688 2472 -2493
rect -2472 -2924 2216 -2688
rect 2452 -2924 2472 -2688
rect -2472 -3008 2472 -2924
rect -2472 -3244 2216 -3008
rect 2452 -3244 2472 -3008
rect -2472 -3328 2472 -3244
rect -2472 -3564 2216 -3328
rect 2452 -3564 2472 -3328
rect -2472 -3648 2472 -3564
rect -2472 -3884 2216 -3648
rect 2452 -3884 2472 -3648
rect -2472 -3968 2472 -3884
rect -2472 -4204 2216 -3968
rect 2452 -4204 2472 -3968
rect -2472 -4288 2472 -4204
rect -2472 -4524 2216 -4288
rect 2452 -4524 2472 -4288
rect -2472 -4608 2472 -4524
rect -2472 -4844 2216 -4608
rect 2452 -4844 2472 -4608
rect -2472 -4928 2472 -4844
rect -2472 -5164 2216 -4928
rect 2452 -5164 2472 -4928
rect -2472 -5248 2472 -5164
rect -2472 -5484 2216 -5248
rect 2452 -5484 2472 -5248
rect -2472 -5568 2472 -5484
rect -2472 -5804 2216 -5568
rect 2452 -5804 2472 -5568
rect -2472 -5888 2472 -5804
rect -2472 -6124 2216 -5888
rect 2452 -6124 2472 -5888
rect -2472 -6208 2472 -6124
rect -2472 -6444 2216 -6208
rect 2452 -6444 2472 -6208
rect -2472 -6528 2472 -6444
rect -2472 -6764 2216 -6528
rect 2452 -6764 2472 -6528
rect -2472 -6848 2472 -6764
rect -2472 -7084 2216 -6848
rect 2452 -7084 2472 -6848
rect -2472 -7279 2472 -7084
<< via4 >>
rect 2216 6848 2452 7084
rect 2216 6528 2452 6764
rect 2216 6208 2452 6444
rect 2216 5888 2452 6124
rect 2216 5568 2452 5804
rect 2216 5248 2452 5484
rect 2216 4928 2452 5164
rect 2216 4608 2452 4844
rect 2216 4288 2452 4524
rect 2216 3968 2452 4204
rect 2216 3648 2452 3884
rect 2216 3328 2452 3564
rect 2216 3008 2452 3244
rect 2216 2688 2452 2924
rect 2216 1962 2452 2198
rect 2216 1642 2452 1878
rect 2216 1322 2452 1558
rect 2216 1002 2452 1238
rect 2216 682 2452 918
rect 2216 362 2452 598
rect 2216 42 2452 278
rect 2216 -278 2452 -42
rect 2216 -598 2452 -362
rect 2216 -918 2452 -682
rect 2216 -1238 2452 -1002
rect 2216 -1558 2452 -1322
rect 2216 -1878 2452 -1642
rect 2216 -2198 2452 -1962
rect 2216 -2924 2452 -2688
rect 2216 -3244 2452 -3008
rect 2216 -3564 2452 -3328
rect 2216 -3884 2452 -3648
rect 2216 -4204 2452 -3968
rect 2216 -4524 2452 -4288
rect 2216 -4844 2452 -4608
rect 2216 -5164 2452 -4928
rect 2216 -5484 2452 -5248
rect 2216 -5804 2452 -5568
rect 2216 -6124 2452 -5888
rect 2216 -6444 2452 -6208
rect 2216 -6764 2452 -6528
rect 2216 -7084 2452 -6848
<< mimcap2 >>
rect -2372 7084 2214 7179
rect -2372 2688 -1797 7084
rect 1639 2688 2214 7084
rect -2372 2593 2214 2688
rect -2372 2198 2214 2293
rect -2372 -2198 -1797 2198
rect 1639 -2198 2214 2198
rect -2372 -2293 2214 -2198
rect -2372 -2688 2214 -2593
rect -2372 -7084 -1797 -2688
rect 1639 -7084 2214 -2688
rect -2372 -7179 2214 -7084
<< mimcap2contact >>
rect -1797 2688 1639 7084
rect -1797 -2198 1639 2198
rect -1797 -7084 1639 -2688
<< metal5 >>
rect -239 7163 81 7329
rect -1905 7084 1747 7163
rect -1905 2688 -1797 7084
rect 1639 2688 1747 7084
rect -1905 2609 1747 2688
rect 2174 7084 2494 7329
rect 2174 6848 2216 7084
rect 2452 6848 2494 7084
rect 2174 6764 2494 6848
rect 2174 6528 2216 6764
rect 2452 6528 2494 6764
rect 2174 6444 2494 6528
rect 2174 6208 2216 6444
rect 2452 6208 2494 6444
rect 2174 6124 2494 6208
rect 2174 5888 2216 6124
rect 2452 5888 2494 6124
rect 2174 5804 2494 5888
rect 2174 5568 2216 5804
rect 2452 5568 2494 5804
rect 2174 5484 2494 5568
rect 2174 5248 2216 5484
rect 2452 5248 2494 5484
rect 2174 5164 2494 5248
rect 2174 4928 2216 5164
rect 2452 4928 2494 5164
rect 2174 4844 2494 4928
rect 2174 4608 2216 4844
rect 2452 4608 2494 4844
rect 2174 4524 2494 4608
rect 2174 4288 2216 4524
rect 2452 4288 2494 4524
rect 2174 4204 2494 4288
rect 2174 3968 2216 4204
rect 2452 3968 2494 4204
rect 2174 3884 2494 3968
rect 2174 3648 2216 3884
rect 2452 3648 2494 3884
rect 2174 3564 2494 3648
rect 2174 3328 2216 3564
rect 2452 3328 2494 3564
rect 2174 3244 2494 3328
rect 2174 3008 2216 3244
rect 2452 3008 2494 3244
rect 2174 2924 2494 3008
rect 2174 2688 2216 2924
rect 2452 2688 2494 2924
rect -239 2277 81 2609
rect -1905 2198 1747 2277
rect -1905 -2198 -1797 2198
rect 1639 -2198 1747 2198
rect -1905 -2277 1747 -2198
rect 2174 2198 2494 2688
rect 2174 1962 2216 2198
rect 2452 1962 2494 2198
rect 2174 1878 2494 1962
rect 2174 1642 2216 1878
rect 2452 1642 2494 1878
rect 2174 1558 2494 1642
rect 2174 1322 2216 1558
rect 2452 1322 2494 1558
rect 2174 1238 2494 1322
rect 2174 1002 2216 1238
rect 2452 1002 2494 1238
rect 2174 918 2494 1002
rect 2174 682 2216 918
rect 2452 682 2494 918
rect 2174 598 2494 682
rect 2174 362 2216 598
rect 2452 362 2494 598
rect 2174 278 2494 362
rect 2174 42 2216 278
rect 2452 42 2494 278
rect 2174 -42 2494 42
rect 2174 -278 2216 -42
rect 2452 -278 2494 -42
rect 2174 -362 2494 -278
rect 2174 -598 2216 -362
rect 2452 -598 2494 -362
rect 2174 -682 2494 -598
rect 2174 -918 2216 -682
rect 2452 -918 2494 -682
rect 2174 -1002 2494 -918
rect 2174 -1238 2216 -1002
rect 2452 -1238 2494 -1002
rect 2174 -1322 2494 -1238
rect 2174 -1558 2216 -1322
rect 2452 -1558 2494 -1322
rect 2174 -1642 2494 -1558
rect 2174 -1878 2216 -1642
rect 2452 -1878 2494 -1642
rect 2174 -1962 2494 -1878
rect 2174 -2198 2216 -1962
rect 2452 -2198 2494 -1962
rect -239 -2609 81 -2277
rect -1905 -2688 1747 -2609
rect -1905 -7084 -1797 -2688
rect 1639 -7084 1747 -2688
rect -1905 -7163 1747 -7084
rect 2174 -2688 2494 -2198
rect 2174 -2924 2216 -2688
rect 2452 -2924 2494 -2688
rect 2174 -3008 2494 -2924
rect 2174 -3244 2216 -3008
rect 2452 -3244 2494 -3008
rect 2174 -3328 2494 -3244
rect 2174 -3564 2216 -3328
rect 2452 -3564 2494 -3328
rect 2174 -3648 2494 -3564
rect 2174 -3884 2216 -3648
rect 2452 -3884 2494 -3648
rect 2174 -3968 2494 -3884
rect 2174 -4204 2216 -3968
rect 2452 -4204 2494 -3968
rect 2174 -4288 2494 -4204
rect 2174 -4524 2216 -4288
rect 2452 -4524 2494 -4288
rect 2174 -4608 2494 -4524
rect 2174 -4844 2216 -4608
rect 2452 -4844 2494 -4608
rect 2174 -4928 2494 -4844
rect 2174 -5164 2216 -4928
rect 2452 -5164 2494 -4928
rect 2174 -5248 2494 -5164
rect 2174 -5484 2216 -5248
rect 2452 -5484 2494 -5248
rect 2174 -5568 2494 -5484
rect 2174 -5804 2216 -5568
rect 2452 -5804 2494 -5568
rect 2174 -5888 2494 -5804
rect 2174 -6124 2216 -5888
rect 2452 -6124 2494 -5888
rect 2174 -6208 2494 -6124
rect 2174 -6444 2216 -6208
rect 2452 -6444 2494 -6208
rect 2174 -6528 2494 -6444
rect 2174 -6764 2216 -6528
rect 2452 -6764 2494 -6528
rect 2174 -6848 2494 -6764
rect 2174 -7084 2216 -6848
rect 2452 -7084 2494 -6848
rect -239 -7329 81 -7163
rect 2174 -7329 2494 -7084
<< properties >>
string FIXED_BBOX -2472 2493 2314 7279
<< end >>
