magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< pwell >>
rect 406174 552950 408226 555450
<< mvpsubdiff >>
rect 406200 555373 408200 555424
rect 406200 553027 406231 555373
rect 408169 553027 408200 555373
rect 406200 552976 408200 553027
<< mvpsubdiffcont >>
rect 406231 553027 408169 555373
<< locali >>
rect 406200 555373 408200 555416
rect 406200 555369 406231 555373
rect 408169 555369 408200 555373
rect 406200 553031 406211 555369
rect 408189 553031 408200 555369
rect 406200 553027 406231 553031
rect 408169 553027 408200 553031
rect 406200 552984 408200 553027
<< viali >>
rect 406211 553031 406231 555369
rect 406231 553031 408169 555369
rect 408169 553031 408189 555369
<< metal1 >>
rect 404800 576600 417600 576800
rect 404800 576598 417610 576600
rect 404800 575202 411206 576598
rect 417594 575202 417610 576598
rect 404800 575200 417610 575202
rect 404800 575000 417600 575200
rect 404800 557786 413600 558000
rect 404800 555814 410402 557786
rect 413398 555814 413600 557786
rect 404800 555600 413600 555814
rect 406000 555369 408400 555600
rect 406000 553031 406211 555369
rect 408189 553031 408400 555369
rect 406000 552800 408400 553031
rect 404800 531382 412600 531600
rect 404800 529218 409826 531382
rect 412374 529218 412600 531382
rect 404800 529000 412600 529218
<< via1 >>
rect 411206 575202 417594 576598
rect 410402 555814 413398 557786
rect 409826 529218 412374 531382
<< metal2 >>
rect 411000 576598 417800 576800
rect 411000 575202 411206 576598
rect 417594 575202 417800 576598
rect 411000 575000 417800 575202
rect 408000 557788 413600 558000
rect 408000 557786 410432 557788
rect 413368 557786 413600 557788
rect 408000 555814 410402 557786
rect 413398 555814 413600 557786
rect 408000 555812 410432 555814
rect 413368 555812 413600 555814
rect 408000 555600 413600 555812
rect 409600 531382 412600 531600
rect 409600 529218 409826 531382
rect 412374 529218 412600 531382
rect 409600 529000 412600 529218
<< via2 >>
rect 411212 575232 417588 576568
rect 410432 557786 413368 557788
rect 410432 555814 413368 557786
rect 410432 555812 413368 555814
rect 409832 529232 412368 531368
<< metal3 >>
rect 411000 576572 417800 576800
rect 411000 575228 411208 576572
rect 417592 575228 417800 576572
rect 411000 575000 417800 575228
rect 408000 557792 413600 558000
rect 408000 555808 410428 557792
rect 413372 555808 413600 557792
rect 408000 555600 413600 555808
rect 409600 531372 412600 531600
rect 409600 529228 409828 531372
rect 412372 529228 412600 531372
rect 409600 529000 412600 529228
<< via3 >>
rect 411208 576568 417592 576572
rect 411208 575232 411212 576568
rect 411212 575232 417588 576568
rect 417588 575232 417592 576568
rect 411208 575228 417592 575232
rect 410428 557788 413372 557792
rect 410428 555812 410432 557788
rect 410432 555812 413368 557788
rect 413368 555812 413372 557788
rect 410428 555808 413372 555812
rect 409828 531368 412372 531372
rect 409828 529232 409832 531368
rect 409832 529232 412368 531368
rect 412368 529232 412372 531368
rect 409828 529228 412372 529232
<< metal4 >>
rect 411000 576572 417800 576800
rect 411000 575228 411208 576572
rect 417592 575228 417800 576572
rect 411000 575000 417800 575228
rect 414200 568980 419160 569360
rect 420000 568980 424960 569360
rect 425800 568980 430760 569360
rect 414200 564080 419160 564460
rect 420000 564080 424960 564460
rect 425800 564100 430760 564480
rect 415600 558000 418600 562200
rect 421200 558000 424200 562200
rect 426600 558000 429600 562200
rect 408000 557792 429600 558000
rect 408000 555808 410428 557792
rect 413372 555808 429600 557792
rect 448160 558768 449820 558800
rect 448160 557252 448232 558768
rect 449748 557252 449820 558768
rect 448160 557220 449820 557252
rect 408000 555600 429600 555808
rect 410200 552600 413200 555600
rect 415600 552000 418600 555600
rect 421200 551800 424200 555600
rect 426600 552400 429600 555600
rect 408600 549540 413780 549920
rect 414200 549540 419380 549920
rect 420200 549560 425380 549940
rect 426000 549560 431180 549940
rect 408600 544440 413780 544820
rect 414200 544440 419380 544820
rect 420200 544440 425380 544820
rect 426000 544440 431180 544820
rect 408600 539320 413780 539700
rect 414200 539320 419380 539700
rect 420200 539320 425380 539700
rect 426000 539320 431180 539700
rect 409600 531378 412600 531600
rect 409600 531372 409862 531378
rect 412338 531372 412600 531378
rect 409600 529228 409828 531372
rect 412372 529228 412600 531372
rect 409600 529222 409862 529228
rect 412338 529222 412600 529228
rect 409600 529000 412600 529222
<< via4 >>
rect 411242 575302 417558 576498
rect 448232 557252 449748 558768
rect 409862 531372 412338 531378
rect 409862 529228 412338 531372
rect 409862 529222 412338 529228
<< metal5 >>
rect 411000 576498 433250 576800
rect 411000 575302 411242 576498
rect 417558 575302 433250 576498
rect 411000 575000 433250 575302
rect 415975 574975 433250 575000
rect 415975 573175 417625 574975
rect 421600 573200 423250 574975
rect 427200 573200 428850 574975
rect 431600 571500 433250 574975
rect 431600 571180 433220 571200
rect 433240 571180 433250 571190
rect 431600 563200 433250 571180
rect 448168 558804 449820 558820
rect 448156 558768 449824 558804
rect 448156 557252 448232 558768
rect 449748 557252 449824 558768
rect 448156 557216 449824 557252
rect 410400 533425 412800 536000
rect 415600 533425 418600 536000
rect 421400 533425 424400 536000
rect 427000 533425 430000 536400
rect 448168 533800 449818 557216
rect 448168 533425 449800 533800
rect 410400 531800 449800 533425
rect 410400 531600 412600 531800
rect 436400 531775 447400 531800
rect 409600 531378 412600 531600
rect 409600 529222 409862 531378
rect 412338 529222 412600 531378
rect 409600 529000 412600 529222
<< rm5 >>
rect 431600 571200 433250 571500
rect 433220 571190 433250 571200
rect 433220 571180 433240 571190
use l0_1  l0_1_0
timestamp 1647143569
transform 1 0 388400 0 1 505600
box 43200 43200 60788 59200
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_0
timestamp 1647143569
transform 1 0 416672 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_1
timestamp 1647143569
transform 1 0 422472 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_4GE4YE  sky130_fd_pr__cap_mim_m3_2_4GE4YE_2
timestamp 1647143569
transform 1 0 428272 0 1 566721
box -2472 -7329 2494 7329
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_0
timestamp 1647143569
transform 1 0 411186 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_1
timestamp 1647143569
transform 1 0 416786 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_2
timestamp 1647143569
transform 1 0 422786 0 1 544626
box -2586 -10228 2608 10228
use sky130_fd_pr__cap_mim_m3_2_8BWDGQ  sky130_fd_pr__cap_mim_m3_2_8BWDGQ_3
timestamp 1647143569
transform 1 0 428586 0 1 544626
box -2586 -10228 2608 10228
<< labels >>
flabel metal1 s 404800 556000 406600 557800 0 FreeSans 2000 0 0 0 gnd
port 1 nsew
flabel metal1 s 404800 529000 407200 531600 0 FreeSans 2000 0 0 0 out
port 2 nsew
flabel metal1 s 404800 575000 406600 576800 0 FreeSans 2000 0 0 0 in
port 3 nsew
<< end >>
