magic
tech sky130A
magscale 1 2
timestamp 1646578768
<< checkpaint >>
rect -4732 -4732 588732 708732
<< pwell >>
rect 345714 628229 371128 629058
<< mvpsubdiff >>
rect 345740 629000 371102 629032
rect 345740 628286 345790 629000
rect 371052 628286 371102 629000
rect 345740 628255 371102 628286
<< mvpsubdiffcont >>
rect 345790 628286 371052 629000
<< locali >>
rect 345748 629000 371094 629032
rect 345748 628286 345790 629000
rect 371052 628286 371094 629000
rect 345748 628255 371094 628286
<< viali >>
rect 357600 628309 359290 628991
<< metal1 >>
rect 357470 629394 359442 629457
rect 357470 628062 357541 629394
rect 359385 628062 359442 629394
rect 357470 627990 359442 628062
<< via1 >>
rect 357541 628991 359385 629394
rect 357541 628309 357600 628991
rect 357600 628309 359290 628991
rect 359290 628309 359385 628991
rect 357541 628062 359385 628309
<< metal2 >>
rect 357470 629396 359442 629457
rect 357470 629394 357555 629396
rect 359371 629394 359442 629396
rect 357470 628062 357541 629394
rect 359385 628062 359442 629394
rect 357470 628060 357555 628062
rect 359371 628060 359442 628062
rect 357470 627990 359442 628060
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 357555 629394 359371 629396
rect 357555 628062 359371 629394
rect 357555 628060 359371 628062
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 700788 173094 704800
rect 170894 690577 173094 700738
rect -800 680242 1700 685242
rect 170894 684353 170922 690577
rect 173066 684353 173094 690577
rect 170894 683764 173094 684353
rect 173394 700786 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 173394 690577 175594 700736
rect 173394 684353 173422 690577
rect 175566 684353 175594 690577
rect 173394 683764 175594 684353
rect 222594 700836 224794 704800
rect 222594 690610 224794 700786
rect 222594 684386 222622 690610
rect 224766 684386 224794 690610
rect 222594 683913 224794 684386
rect 225094 700846 227294 704800
rect 227594 702300 232594 704800
rect 225094 690610 227294 700796
rect 225094 684386 225122 690610
rect 227266 684386 227294 690610
rect 225094 683913 227294 684386
rect 318994 649490 323994 704800
rect 324294 701130 326494 704800
rect 324294 690593 326494 701080
rect 326794 701150 328994 704800
rect 326794 694292 328994 701100
rect 329294 694292 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 326794 692092 334294 694292
rect 324294 684369 324322 690593
rect 326466 684369 326494 690593
rect 324294 684038 326494 684369
rect -800 643842 1660 648642
rect 318994 643746 319022 649490
rect 323966 643746 323994 649490
rect 318994 642983 323994 643746
rect 329294 649490 334294 692092
rect 329294 643746 329322 649490
rect 334266 643746 334294 649490
rect 329294 642983 334294 643746
rect 510594 690560 515394 704800
rect 510594 684336 510602 690560
rect 515386 684336 515394 690560
rect -800 633842 1660 638642
rect 510594 637561 515394 684336
rect 510594 631817 510602 637561
rect 515386 631817 515394 637561
rect 510594 631116 515394 631817
rect 520594 690560 525394 704800
rect 566594 702300 571594 704800
rect 520594 684336 520602 690560
rect 525386 684336 525394 690560
rect 520594 637561 525394 684336
rect 582300 677984 584800 682984
rect 560050 644576 584800 644584
rect 560050 639792 560582 644576
rect 566726 639792 584800 644576
rect 560050 639784 584800 639792
rect 520594 631817 520602 637561
rect 525386 631817 525394 637561
rect 520594 631116 525394 631817
rect 560050 634576 584800 634584
rect 560050 629792 560582 634576
rect 566726 629792 584800 634576
rect 560050 629784 584800 629792
rect 357470 629396 359442 629457
rect 357470 629360 357555 629396
rect 359371 629360 359442 629396
rect 357470 628096 357551 629360
rect 359375 628096 359442 629360
rect 357470 628060 357555 628096
rect 359371 628060 359442 628096
rect 357470 627990 359442 628060
rect 339960 620294 345660 620363
rect 371099 620302 533609 620371
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 339960 511642 340072 620294
rect 341733 619661 341855 619684
rect 341733 619597 341762 619661
rect 341826 619637 341855 619661
rect 533089 619645 533095 619647
rect 341826 619597 345660 619637
rect 341733 619577 345660 619597
rect 371099 619585 533095 619645
rect 533089 619583 533095 619585
rect 533159 619583 533165 619647
rect 341733 619574 341855 619577
rect 533105 619280 533111 619282
rect -800 511530 340072 511642
rect 340967 619212 345660 619272
rect 371099 619220 533111 619280
rect 533105 619218 533111 619220
rect 533175 619218 533181 619282
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect 340967 463692 341079 619212
rect -800 463580 341079 463692
rect 341738 618608 341850 618638
rect 341738 618544 341762 618608
rect 341826 618544 341850 618608
rect -800 462398 660 462510
rect 780 462486 17711 462510
rect 780 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17711 462486
rect 780 462398 17711 462422
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 341738 420470 341850 618544
rect -800 420358 341850 420470
rect -800 419176 676 419288
rect 738 419264 17694 419288
rect 738 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17694 419264
rect 738 419176 17694 419200
rect 533497 405408 533609 620302
rect 533894 619647 533958 619653
rect 533958 619585 539606 619645
rect 533894 619577 533958 619583
rect 533904 619282 533968 619288
rect 533968 619220 537488 619280
rect 533904 619212 533968 619218
rect 537376 454558 537488 619220
rect 539494 498980 539606 619585
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 555452 555354 584800 555362
rect 555452 550570 556255 555354
rect 562319 550570 584800 555354
rect 555452 550562 584800 550570
rect 555452 545354 584800 545362
rect 555452 540570 556255 545354
rect 562319 540570 584800 545354
rect 555452 540562 584800 540570
rect 573371 500138 583220 500162
rect 573371 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 583220 500138
rect 573371 500050 583220 500074
rect 583318 500050 584800 500162
rect 539494 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 573405 455716 583180 455740
rect 573405 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 583180 455716
rect 573405 455628 583180 455652
rect 583296 455628 584800 455740
rect 537376 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 533497 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 13406 196222 584800 196230
rect 13406 191438 13997 196222
rect 17421 191438 573605 196222
rect 576629 191438 584800 196222
rect 13406 191430 584800 191438
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< rmetal3 >>
rect 170894 700738 173094 700788
rect 173394 700736 175594 700786
rect 222594 700786 224794 700836
rect 225094 700796 227294 700846
rect 324294 701080 326494 701130
rect 326794 701100 328994 701150
rect 660 462398 780 462510
rect 676 419176 738 419288
rect 583220 500050 583318 500162
rect 583180 455628 583296 455740
<< via3 >>
rect 170922 684353 173066 690577
rect 173422 684353 175566 690577
rect 222622 684386 224766 690610
rect 225122 684386 227266 690610
rect 324322 684369 326466 690593
rect 319022 643746 323966 649490
rect 329322 643746 334266 649490
rect 510602 684336 515386 690560
rect 510602 631817 515386 637561
rect 520602 684336 525386 690560
rect 560582 639792 566726 644576
rect 520602 631817 525386 637561
rect 560582 629792 566726 634576
rect 357551 628096 357555 629360
rect 357555 628096 359371 629360
rect 359371 628096 359375 629360
rect 341762 619597 341826 619661
rect 533095 619583 533159 619647
rect 533111 619218 533175 619282
rect 341762 618544 341826 618608
rect 13897 462422 13961 462486
rect 13977 462422 14041 462486
rect 14057 462422 14121 462486
rect 14137 462422 14201 462486
rect 14217 462422 14281 462486
rect 14297 462422 14361 462486
rect 14377 462422 14441 462486
rect 14457 462422 14521 462486
rect 14537 462422 14601 462486
rect 14617 462422 14681 462486
rect 14697 462422 14761 462486
rect 14777 462422 14841 462486
rect 14857 462422 14921 462486
rect 14937 462422 15001 462486
rect 15017 462422 15081 462486
rect 15097 462422 15161 462486
rect 15177 462422 15241 462486
rect 15257 462422 15321 462486
rect 15337 462422 15401 462486
rect 15417 462422 15481 462486
rect 15497 462422 15561 462486
rect 15577 462422 15641 462486
rect 15657 462422 15721 462486
rect 15737 462422 15801 462486
rect 15817 462422 15881 462486
rect 15897 462422 15961 462486
rect 15977 462422 16041 462486
rect 16057 462422 16121 462486
rect 16137 462422 16201 462486
rect 16217 462422 16281 462486
rect 16297 462422 16361 462486
rect 16377 462422 16441 462486
rect 16457 462422 16521 462486
rect 16537 462422 16601 462486
rect 16617 462422 16681 462486
rect 16697 462422 16761 462486
rect 16777 462422 16841 462486
rect 16857 462422 16921 462486
rect 16937 462422 17001 462486
rect 17017 462422 17081 462486
rect 17097 462422 17161 462486
rect 17177 462422 17241 462486
rect 17257 462422 17321 462486
rect 17337 462422 17401 462486
rect 17417 462422 17481 462486
rect 17497 462422 17561 462486
rect 13911 419200 13975 419264
rect 13991 419200 14055 419264
rect 14071 419200 14135 419264
rect 14151 419200 14215 419264
rect 14231 419200 14295 419264
rect 14311 419200 14375 419264
rect 14391 419200 14455 419264
rect 14471 419200 14535 419264
rect 14551 419200 14615 419264
rect 14631 419200 14695 419264
rect 14711 419200 14775 419264
rect 14791 419200 14855 419264
rect 14871 419200 14935 419264
rect 14951 419200 15015 419264
rect 15031 419200 15095 419264
rect 15111 419200 15175 419264
rect 15191 419200 15255 419264
rect 15271 419200 15335 419264
rect 15351 419200 15415 419264
rect 15431 419200 15495 419264
rect 15511 419200 15575 419264
rect 15591 419200 15655 419264
rect 15671 419200 15735 419264
rect 15751 419200 15815 419264
rect 15831 419200 15895 419264
rect 15911 419200 15975 419264
rect 15991 419200 16055 419264
rect 16071 419200 16135 419264
rect 16151 419200 16215 419264
rect 16231 419200 16295 419264
rect 16311 419200 16375 419264
rect 16391 419200 16455 419264
rect 16471 419200 16535 419264
rect 16551 419200 16615 419264
rect 16631 419200 16695 419264
rect 16711 419200 16775 419264
rect 16791 419200 16855 419264
rect 16871 419200 16935 419264
rect 16951 419200 17015 419264
rect 17031 419200 17095 419264
rect 17111 419200 17175 419264
rect 17191 419200 17255 419264
rect 17271 419200 17335 419264
rect 17351 419200 17415 419264
rect 17431 419200 17495 419264
rect 17511 419200 17575 419264
rect 533894 619583 533958 619647
rect 533904 619218 533968 619282
rect 556255 550570 562319 555354
rect 556255 540570 562319 545354
rect 573553 500074 573617 500138
rect 573633 500074 573697 500138
rect 573713 500074 573777 500138
rect 573793 500074 573857 500138
rect 573873 500074 573937 500138
rect 573953 500074 574017 500138
rect 574033 500074 574097 500138
rect 574113 500074 574177 500138
rect 574193 500074 574257 500138
rect 574273 500074 574337 500138
rect 574353 500074 574417 500138
rect 574433 500074 574497 500138
rect 574513 500074 574577 500138
rect 574593 500074 574657 500138
rect 574673 500074 574737 500138
rect 574753 500074 574817 500138
rect 574833 500074 574897 500138
rect 574913 500074 574977 500138
rect 574993 500074 575057 500138
rect 575073 500074 575137 500138
rect 575153 500074 575217 500138
rect 575233 500074 575297 500138
rect 575313 500074 575377 500138
rect 575393 500074 575457 500138
rect 575473 500074 575537 500138
rect 575553 500074 575617 500138
rect 575633 500074 575697 500138
rect 575713 500074 575777 500138
rect 575793 500074 575857 500138
rect 575873 500074 575937 500138
rect 575953 500074 576017 500138
rect 576033 500074 576097 500138
rect 576113 500074 576177 500138
rect 576193 500074 576257 500138
rect 576273 500074 576337 500138
rect 576353 500074 576417 500138
rect 576433 500074 576497 500138
rect 576513 500074 576577 500138
rect 576593 500074 576657 500138
rect 576673 500074 576737 500138
rect 573591 455652 573655 455716
rect 573671 455652 573735 455716
rect 573751 455652 573815 455716
rect 573831 455652 573895 455716
rect 573911 455652 573975 455716
rect 573991 455652 574055 455716
rect 574071 455652 574135 455716
rect 574151 455652 574215 455716
rect 574231 455652 574295 455716
rect 574311 455652 574375 455716
rect 574391 455652 574455 455716
rect 574471 455652 574535 455716
rect 574551 455652 574615 455716
rect 574631 455652 574695 455716
rect 574711 455652 574775 455716
rect 574791 455652 574855 455716
rect 574871 455652 574935 455716
rect 574951 455652 575015 455716
rect 575031 455652 575095 455716
rect 575111 455652 575175 455716
rect 575191 455652 575255 455716
rect 575271 455652 575335 455716
rect 575351 455652 575415 455716
rect 575431 455652 575495 455716
rect 575511 455652 575575 455716
rect 575591 455652 575655 455716
rect 575671 455652 575735 455716
rect 575751 455652 575815 455716
rect 575831 455652 575895 455716
rect 575911 455652 575975 455716
rect 575991 455652 576055 455716
rect 576071 455652 576135 455716
rect 576151 455652 576215 455716
rect 576231 455652 576295 455716
rect 576311 455652 576375 455716
rect 576391 455652 576455 455716
rect 576471 455652 576535 455716
rect 576551 455652 576615 455716
rect 576631 455652 576695 455716
rect 13997 191438 17421 196222
rect 573605 191438 576629 196222
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 170628 690610 526162 690737
rect 170628 690577 222622 690610
rect 170628 684353 170922 690577
rect 173066 684353 173422 690577
rect 175566 684386 222622 690577
rect 224766 684386 225122 690610
rect 227266 690593 526162 690610
rect 227266 684386 324322 690593
rect 175566 684369 324322 684386
rect 326466 690560 526162 690593
rect 326466 684369 510602 690560
rect 175566 684353 510602 684369
rect 170628 684336 510602 684353
rect 515386 684336 520602 690560
rect 525386 684336 526162 690560
rect 170628 684183 526162 684336
rect 318330 649773 359973 649898
rect 318330 649490 357678 649773
rect 318330 643746 319022 649490
rect 323966 643746 329322 649490
rect 334266 643746 357678 649490
rect 318330 643457 357678 643746
rect 359194 643457 359973 649773
rect 318330 643344 359973 643457
rect 560425 644576 566979 644980
rect 560425 639792 560582 644576
rect 566726 639792 566979 644576
rect 356144 637561 525696 637898
rect 356144 631817 510602 637561
rect 515386 631817 520602 637561
rect 525386 631817 525696 637561
rect 356144 631344 525696 631817
rect 560425 634576 566979 639792
rect 357442 629360 359470 631344
rect 357442 628096 357551 629360
rect 359375 628096 359470 629360
rect 357442 619873 359470 628096
rect 560425 629792 560582 634576
rect 566726 629792 566979 634576
rect 341738 619661 341850 619685
rect 341738 619597 341762 619661
rect 341826 619597 341850 619661
rect 341738 618633 341850 619597
rect 356867 619473 359885 619873
rect 533094 619647 533160 619648
rect 533094 619583 533095 619647
rect 533159 619645 533160 619647
rect 533893 619647 533959 619648
rect 533893 619645 533894 619647
rect 533159 619585 533894 619645
rect 533159 619583 533160 619585
rect 533094 619582 533160 619583
rect 533893 619583 533894 619585
rect 533958 619583 533959 619647
rect 533893 619582 533959 619583
rect 533110 619282 533176 619283
rect 533110 619218 533111 619282
rect 533175 619280 533176 619282
rect 533903 619282 533969 619283
rect 533903 619280 533904 619282
rect 533175 619220 533904 619280
rect 533175 619218 533176 619220
rect 533110 619217 533176 619218
rect 533903 619218 533904 619220
rect 533968 619218 533969 619282
rect 533903 619217 533969 619218
rect 341737 618608 341851 618633
rect 341737 618544 341762 618608
rect 341826 618544 341851 618608
rect 341737 618519 341851 618544
rect 345773 613756 346828 618849
rect 351928 617777 353757 618856
rect 351928 615301 352057 617777
rect 353573 615301 353757 617777
rect 351928 615131 353757 615301
rect 363328 617783 365157 618884
rect 363328 615307 363441 617783
rect 364957 615307 365157 617783
rect 363328 615131 365157 615307
rect 369823 613756 370980 618859
rect 560425 613756 566979 629792
rect 345256 607202 566979 613756
rect 362658 601439 562613 601756
rect 362658 597363 363445 601439
rect 364961 597363 562613 601439
rect 362658 595202 562613 597363
rect 556059 555354 562613 595202
rect 556059 550570 556255 555354
rect 562319 550570 562613 555354
rect 556059 545354 562613 550570
rect 556059 540570 556255 545354
rect 562319 540570 562613 545354
rect 556059 540155 562613 540570
rect 573464 500138 576816 500473
rect 573464 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 576816 500138
rect 13814 462486 17684 462771
rect 13814 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17684 462486
rect 13814 419264 17684 462422
rect 13814 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17684 419264
rect 13814 227257 17684 419200
rect 573464 455716 576816 500074
rect 573464 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 576816 455716
rect 13811 196222 17688 227257
rect 13811 191438 13997 196222
rect 17421 191438 17688 196222
rect 13811 191098 17688 191438
rect 573464 196222 576816 455652
rect 573464 191438 573605 196222
rect 576629 191438 576816 196222
rect 573464 191191 576816 191438
<< via4 >>
rect 357678 643457 359194 649773
rect 352057 615301 353573 617777
rect 363441 615307 364957 617783
rect 363445 597363 364961 601439
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 357521 649773 359350 649991
rect 357521 643457 357678 649773
rect 359194 643457 359350 649773
rect 351918 617777 353747 617929
rect 351918 615301 352057 617777
rect 353573 615301 353747 617777
rect 351918 614900 353747 615301
rect 357521 614900 359350 643457
rect 351918 613071 359350 614900
rect 363318 617783 365147 617929
rect 363318 615307 363441 617783
rect 364957 615307 365147 617783
rect 363318 601439 365147 615307
rect 363318 597363 363445 601439
rect 364961 597363 365147 601439
rect 363318 597052 365147 597363
use user_analog_proj_example  user_analog_proj_example_0
timestamp 1639823760
transform 1 0 345668 0 -1 627114
box -73 -12 25490 8324
<< labels >>
flabel metal3 s 572152 640142 580220 644150 0 FreeSans 20000 0 0 0 VCCD1
port 1 nsew
flabel metal3 s 567038 550960 577302 554546 0 FreeSans 20000 0 0 0 VDDA1
port 2 nsew
flabel metal3 s 511190 664896 514962 676272 0 FreeSans 20000 90 0 0 VSSA1
port 3 nsew
flabel metal3 s 561703 191929 571721 195859 0 FreeSans 20000 0 0 0 VSSD1
port 4 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 5 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 6 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 7 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 8 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 9 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 10 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 11 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 12 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 13 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 14 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 15 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 16 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 17 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 18 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 19 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 20 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 21 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 22 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 23 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 24 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 25 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 26 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 27 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 28 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 29 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 30 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 31 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 32 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 33 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 34 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 35 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 36 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 37 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 38 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 39 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 40 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 41 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 42 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 43 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 44 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 45 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 49 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 50 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 51 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 46 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 47 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 48 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 52 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 53 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 54 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 55 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 56 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 57 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 58 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 59 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 60 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 61 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 62 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 63 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 64 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 65 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 66 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 67 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 68 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 69 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 70 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 71 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 72 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 73 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 74 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 75 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 76 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 77 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 78 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 79 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 80 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 81 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 82 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 83 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 84 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 85 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 86 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 87 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 88 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 89 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 90 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 91 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 92 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 93 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 94 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 95 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 96 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 97 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 98 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 99 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 100 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 101 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 102 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 103 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 104 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 105 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 106 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 107 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 108 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 109 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 110 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 111 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 112 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 113 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 114 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 115 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 116 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 117 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 118 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 119 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 120 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 121 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 122 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 123 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 124 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 125 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 126 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 127 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 128 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 129 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 130 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 131 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 132 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 133 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 134 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 135 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 136 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 137 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 138 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 139 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 140 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 141 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 142 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 143 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 144 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 145 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 146 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 147 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 148 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 149 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 150 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 151 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 152 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 153 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 154 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 155 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 156 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 157 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 158 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 159 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 160 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 161 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 162 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 163 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 164 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 165 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 166 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 167 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 168 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 169 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 170 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 171 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 172 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 173 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 174 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 175 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 176 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 177 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 178 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 179 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 180 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 181 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 182 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 183 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 184 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 185 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 186 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 187 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 188 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 189 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 190 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 191 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 192 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 193 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 194 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 195 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 196 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 197 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 198 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 199 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 200 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 201 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 202 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 203 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 204 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 205 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 206 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 207 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 208 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 209 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 210 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 211 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 212 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 213 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 214 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 215 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 216 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 217 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 218 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 219 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 220 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 221 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 222 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 223 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 224 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 225 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 226 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 227 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 228 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 229 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 230 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 231 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 232 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 233 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 234 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 235 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 236 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 237 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 238 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 239 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 240 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 241 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 242 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 243 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 244 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 245 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 246 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 247 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 248 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 249 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 250 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 251 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 252 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 253 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 254 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 255 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 256 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 257 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 258 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 259 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 260 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 261 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 262 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 263 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 264 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 265 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 266 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 267 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 268 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 269 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 270 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 271 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 272 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 273 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 274 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 275 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 276 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 277 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 278 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 279 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 280 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 281 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 282 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 283 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 284 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 285 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 286 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 287 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 288 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 289 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 290 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 291 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 292 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 293 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 294 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 295 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 296 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 297 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 298 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 299 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 300 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 301 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 302 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 303 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 304 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 305 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 306 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 307 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 308 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 309 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 310 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 311 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 312 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 313 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 314 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 315 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 316 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 317 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 318 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 319 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 320 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 321 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 322 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 323 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 324 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 325 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 326 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 327 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 328 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 329 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 330 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 331 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 332 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 333 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 334 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 335 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 336 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 337 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 338 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 339 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 340 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 341 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 342 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 343 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 344 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 345 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 346 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 347 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 348 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 349 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 350 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 351 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 352 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 353 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 354 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 355 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 356 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 357 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 358 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 359 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 360 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 361 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 362 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 363 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 364 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 365 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 366 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 367 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 368 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 369 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 370 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 371 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 372 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 373 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 374 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 375 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 376 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 377 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 378 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 379 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 380 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 381 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 382 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 383 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 384 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 385 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 386 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 387 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 388 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 389 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 390 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 391 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 392 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 393 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 394 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 395 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 396 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 397 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 398 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 399 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 400 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 401 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 402 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 403 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 404 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 405 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 406 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 407 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 408 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 409 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 410 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 411 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 412 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 413 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 414 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 415 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 416 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 417 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 418 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 419 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 420 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 421 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 422 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 423 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 424 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 425 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 426 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 427 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 428 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 429 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 430 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 431 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 432 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 433 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 434 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 435 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 436 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 437 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 438 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 439 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 440 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 441 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 442 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 443 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 444 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 445 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 446 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 447 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 448 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 449 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 450 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 451 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 452 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 453 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 454 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 455 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 456 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 457 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 458 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 459 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 460 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 461 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 462 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 463 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 464 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 465 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 466 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 467 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 468 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 469 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 470 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 471 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 472 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 473 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 474 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 475 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 476 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 477 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 478 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 479 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 480 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 481 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 482 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 483 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 484 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 485 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 486 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 487 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 488 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 489 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 490 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 491 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 492 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 493 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 494 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 495 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 496 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 497 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 498 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 499 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 500 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 501 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 502 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 503 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 504 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 505 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 506 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 507 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 508 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 509 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 510 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 511 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 512 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 513 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 514 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 515 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 516 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 517 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 518 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 519 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 520 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 521 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 522 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 523 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 524 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 525 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 526 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 527 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 528 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 529 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 530 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 531 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 532 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 533 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 534 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 535 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 536 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 537 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 538 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 539 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 540 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 541 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 542 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 543 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 544 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 545 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 546 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 547 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 548 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 549 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 550 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 551 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 552 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 553 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 554 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 554 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 555 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 555 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 556 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 556 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 556 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 556 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 557 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 557 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 558 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 558 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 558 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 558 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 559 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 559 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 560 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 560 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 561 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 561 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 562 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 563 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 564 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 565 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 566 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 567 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 568 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 569 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 570 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 571 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 572 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 573 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 574 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 575 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 576 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 577 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 578 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 579 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 580 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 581 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 582 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 583 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 584 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 585 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 586 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 587 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 588 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 589 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 590 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 591 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 592 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 593 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 594 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 595 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 596 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 597 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 598 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 599 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 600 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 601 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 602 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 603 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 604 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 605 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 606 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 607 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 608 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 609 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 610 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 611 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 612 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 613 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 614 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 615 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 616 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 617 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 618 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 619 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 620 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 621 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 622 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 623 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 624 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 625 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 626 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 627 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 628 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 629 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 630 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 631 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 632 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 633 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 634 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 635 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 636 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 637 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 638 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 639 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 640 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 641 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 642 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 643 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 644 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 645 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 646 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 647 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 648 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 649 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 650 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 651 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 652 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 653 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 654 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 655 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 656 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 657 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 658 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 659 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 660 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 661 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 662 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 663 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 664 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 665 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 666 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 667 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
