magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< metal4 >>
rect -2619 7538 2619 7720
rect -2619 7302 2363 7538
rect 2599 7302 2619 7538
rect -2619 7218 2619 7302
rect -2619 6982 2363 7218
rect 2599 6982 2619 7218
rect -2619 6898 2619 6982
rect -2619 6662 2363 6898
rect 2599 6662 2619 6898
rect -2619 6578 2619 6662
rect -2619 6342 2363 6578
rect 2599 6342 2619 6578
rect -2619 6258 2619 6342
rect -2619 6022 2363 6258
rect 2599 6022 2619 6258
rect -2619 5938 2619 6022
rect -2619 5702 2363 5938
rect 2599 5702 2619 5938
rect -2619 5618 2619 5702
rect -2619 5382 2363 5618
rect 2599 5382 2619 5618
rect -2619 5298 2619 5382
rect -2619 5062 2363 5298
rect 2599 5062 2619 5298
rect -2619 4978 2619 5062
rect -2619 4742 2363 4978
rect 2599 4742 2619 4978
rect -2619 4658 2619 4742
rect -2619 4422 2363 4658
rect 2599 4422 2619 4658
rect -2619 4338 2619 4422
rect -2619 4102 2363 4338
rect 2599 4102 2619 4338
rect -2619 4018 2619 4102
rect -2619 3782 2363 4018
rect 2599 3782 2619 4018
rect -2619 3698 2619 3782
rect -2619 3462 2363 3698
rect 2599 3462 2619 3698
rect -2619 3378 2619 3462
rect -2619 3142 2363 3378
rect 2599 3142 2619 3378
rect -2619 3058 2619 3142
rect -2619 2822 2363 3058
rect 2599 2822 2619 3058
rect -2619 2640 2619 2822
rect -2619 2358 2619 2540
rect -2619 2122 2363 2358
rect 2599 2122 2619 2358
rect -2619 2038 2619 2122
rect -2619 1802 2363 2038
rect 2599 1802 2619 2038
rect -2619 1718 2619 1802
rect -2619 1482 2363 1718
rect 2599 1482 2619 1718
rect -2619 1398 2619 1482
rect -2619 1162 2363 1398
rect 2599 1162 2619 1398
rect -2619 1078 2619 1162
rect -2619 842 2363 1078
rect 2599 842 2619 1078
rect -2619 758 2619 842
rect -2619 522 2363 758
rect 2599 522 2619 758
rect -2619 438 2619 522
rect -2619 202 2363 438
rect 2599 202 2619 438
rect -2619 118 2619 202
rect -2619 -118 2363 118
rect 2599 -118 2619 118
rect -2619 -202 2619 -118
rect -2619 -438 2363 -202
rect 2599 -438 2619 -202
rect -2619 -522 2619 -438
rect -2619 -758 2363 -522
rect 2599 -758 2619 -522
rect -2619 -842 2619 -758
rect -2619 -1078 2363 -842
rect 2599 -1078 2619 -842
rect -2619 -1162 2619 -1078
rect -2619 -1398 2363 -1162
rect 2599 -1398 2619 -1162
rect -2619 -1482 2619 -1398
rect -2619 -1718 2363 -1482
rect 2599 -1718 2619 -1482
rect -2619 -1802 2619 -1718
rect -2619 -2038 2363 -1802
rect 2599 -2038 2619 -1802
rect -2619 -2122 2619 -2038
rect -2619 -2358 2363 -2122
rect 2599 -2358 2619 -2122
rect -2619 -2540 2619 -2358
rect -2619 -2822 2619 -2640
rect -2619 -3058 2363 -2822
rect 2599 -3058 2619 -2822
rect -2619 -3142 2619 -3058
rect -2619 -3378 2363 -3142
rect 2599 -3378 2619 -3142
rect -2619 -3462 2619 -3378
rect -2619 -3698 2363 -3462
rect 2599 -3698 2619 -3462
rect -2619 -3782 2619 -3698
rect -2619 -4018 2363 -3782
rect 2599 -4018 2619 -3782
rect -2619 -4102 2619 -4018
rect -2619 -4338 2363 -4102
rect 2599 -4338 2619 -4102
rect -2619 -4422 2619 -4338
rect -2619 -4658 2363 -4422
rect 2599 -4658 2619 -4422
rect -2619 -4742 2619 -4658
rect -2619 -4978 2363 -4742
rect 2599 -4978 2619 -4742
rect -2619 -5062 2619 -4978
rect -2619 -5298 2363 -5062
rect 2599 -5298 2619 -5062
rect -2619 -5382 2619 -5298
rect -2619 -5618 2363 -5382
rect 2599 -5618 2619 -5382
rect -2619 -5702 2619 -5618
rect -2619 -5938 2363 -5702
rect 2599 -5938 2619 -5702
rect -2619 -6022 2619 -5938
rect -2619 -6258 2363 -6022
rect 2599 -6258 2619 -6022
rect -2619 -6342 2619 -6258
rect -2619 -6578 2363 -6342
rect 2599 -6578 2619 -6342
rect -2619 -6662 2619 -6578
rect -2619 -6898 2363 -6662
rect 2599 -6898 2619 -6662
rect -2619 -6982 2619 -6898
rect -2619 -7218 2363 -6982
rect 2599 -7218 2619 -6982
rect -2619 -7302 2619 -7218
rect -2619 -7538 2363 -7302
rect 2599 -7538 2619 -7302
rect -2619 -7720 2619 -7538
<< via4 >>
rect 2363 7302 2599 7538
rect 2363 6982 2599 7218
rect 2363 6662 2599 6898
rect 2363 6342 2599 6578
rect 2363 6022 2599 6258
rect 2363 5702 2599 5938
rect 2363 5382 2599 5618
rect 2363 5062 2599 5298
rect 2363 4742 2599 4978
rect 2363 4422 2599 4658
rect 2363 4102 2599 4338
rect 2363 3782 2599 4018
rect 2363 3462 2599 3698
rect 2363 3142 2599 3378
rect 2363 2822 2599 3058
rect 2363 2122 2599 2358
rect 2363 1802 2599 2038
rect 2363 1482 2599 1718
rect 2363 1162 2599 1398
rect 2363 842 2599 1078
rect 2363 522 2599 758
rect 2363 202 2599 438
rect 2363 -118 2599 118
rect 2363 -438 2599 -202
rect 2363 -758 2599 -522
rect 2363 -1078 2599 -842
rect 2363 -1398 2599 -1162
rect 2363 -1718 2599 -1482
rect 2363 -2038 2599 -1802
rect 2363 -2358 2599 -2122
rect 2363 -3058 2599 -2822
rect 2363 -3378 2599 -3142
rect 2363 -3698 2599 -3462
rect 2363 -4018 2599 -3782
rect 2363 -4338 2599 -4102
rect 2363 -4658 2599 -4422
rect 2363 -4978 2599 -4742
rect 2363 -5298 2599 -5062
rect 2363 -5618 2599 -5382
rect 2363 -5938 2599 -5702
rect 2363 -6258 2599 -6022
rect 2363 -6578 2599 -6342
rect 2363 -6898 2599 -6662
rect 2363 -7218 2599 -6982
rect 2363 -7538 2599 -7302
<< mimcap2 >>
rect -2519 7538 2361 7620
rect -2519 2822 -1957 7538
rect 1799 2822 2361 7538
rect -2519 2740 2361 2822
rect -2519 2358 2361 2440
rect -2519 -2358 -1957 2358
rect 1799 -2358 2361 2358
rect -2519 -2440 2361 -2358
rect -2519 -2822 2361 -2740
rect -2519 -7538 -1957 -2822
rect 1799 -7538 2361 -2822
rect -2519 -7620 2361 -7538
<< mimcap2contact >>
rect -1957 2822 1799 7538
rect -1957 -2358 1799 2358
rect -1957 -7538 1799 -2822
<< metal5 >>
rect -239 7604 81 7770
rect -2023 7538 1865 7604
rect -2023 2822 -1957 7538
rect 1799 2822 1865 7538
rect -2023 2756 1865 2822
rect 2321 7538 2641 7770
rect 2321 7302 2363 7538
rect 2599 7302 2641 7538
rect 2321 7218 2641 7302
rect 2321 6982 2363 7218
rect 2599 6982 2641 7218
rect 2321 6898 2641 6982
rect 2321 6662 2363 6898
rect 2599 6662 2641 6898
rect 2321 6578 2641 6662
rect 2321 6342 2363 6578
rect 2599 6342 2641 6578
rect 2321 6258 2641 6342
rect 2321 6022 2363 6258
rect 2599 6022 2641 6258
rect 2321 5938 2641 6022
rect 2321 5702 2363 5938
rect 2599 5702 2641 5938
rect 2321 5618 2641 5702
rect 2321 5382 2363 5618
rect 2599 5382 2641 5618
rect 2321 5298 2641 5382
rect 2321 5062 2363 5298
rect 2599 5062 2641 5298
rect 2321 4978 2641 5062
rect 2321 4742 2363 4978
rect 2599 4742 2641 4978
rect 2321 4658 2641 4742
rect 2321 4422 2363 4658
rect 2599 4422 2641 4658
rect 2321 4338 2641 4422
rect 2321 4102 2363 4338
rect 2599 4102 2641 4338
rect 2321 4018 2641 4102
rect 2321 3782 2363 4018
rect 2599 3782 2641 4018
rect 2321 3698 2641 3782
rect 2321 3462 2363 3698
rect 2599 3462 2641 3698
rect 2321 3378 2641 3462
rect 2321 3142 2363 3378
rect 2599 3142 2641 3378
rect 2321 3058 2641 3142
rect 2321 2822 2363 3058
rect 2599 2822 2641 3058
rect -239 2424 81 2756
rect -2023 2358 1865 2424
rect -2023 -2358 -1957 2358
rect 1799 -2358 1865 2358
rect -2023 -2424 1865 -2358
rect 2321 2358 2641 2822
rect 2321 2122 2363 2358
rect 2599 2122 2641 2358
rect 2321 2038 2641 2122
rect 2321 1802 2363 2038
rect 2599 1802 2641 2038
rect 2321 1718 2641 1802
rect 2321 1482 2363 1718
rect 2599 1482 2641 1718
rect 2321 1398 2641 1482
rect 2321 1162 2363 1398
rect 2599 1162 2641 1398
rect 2321 1078 2641 1162
rect 2321 842 2363 1078
rect 2599 842 2641 1078
rect 2321 758 2641 842
rect 2321 522 2363 758
rect 2599 522 2641 758
rect 2321 438 2641 522
rect 2321 202 2363 438
rect 2599 202 2641 438
rect 2321 118 2641 202
rect 2321 -118 2363 118
rect 2599 -118 2641 118
rect 2321 -202 2641 -118
rect 2321 -438 2363 -202
rect 2599 -438 2641 -202
rect 2321 -522 2641 -438
rect 2321 -758 2363 -522
rect 2599 -758 2641 -522
rect 2321 -842 2641 -758
rect 2321 -1078 2363 -842
rect 2599 -1078 2641 -842
rect 2321 -1162 2641 -1078
rect 2321 -1398 2363 -1162
rect 2599 -1398 2641 -1162
rect 2321 -1482 2641 -1398
rect 2321 -1718 2363 -1482
rect 2599 -1718 2641 -1482
rect 2321 -1802 2641 -1718
rect 2321 -2038 2363 -1802
rect 2599 -2038 2641 -1802
rect 2321 -2122 2641 -2038
rect 2321 -2358 2363 -2122
rect 2599 -2358 2641 -2122
rect -239 -2756 81 -2424
rect -2023 -2822 1865 -2756
rect -2023 -7538 -1957 -2822
rect 1799 -7538 1865 -2822
rect -2023 -7604 1865 -7538
rect 2321 -2822 2641 -2358
rect 2321 -3058 2363 -2822
rect 2599 -3058 2641 -2822
rect 2321 -3142 2641 -3058
rect 2321 -3378 2363 -3142
rect 2599 -3378 2641 -3142
rect 2321 -3462 2641 -3378
rect 2321 -3698 2363 -3462
rect 2599 -3698 2641 -3462
rect 2321 -3782 2641 -3698
rect 2321 -4018 2363 -3782
rect 2599 -4018 2641 -3782
rect 2321 -4102 2641 -4018
rect 2321 -4338 2363 -4102
rect 2599 -4338 2641 -4102
rect 2321 -4422 2641 -4338
rect 2321 -4658 2363 -4422
rect 2599 -4658 2641 -4422
rect 2321 -4742 2641 -4658
rect 2321 -4978 2363 -4742
rect 2599 -4978 2641 -4742
rect 2321 -5062 2641 -4978
rect 2321 -5298 2363 -5062
rect 2599 -5298 2641 -5062
rect 2321 -5382 2641 -5298
rect 2321 -5618 2363 -5382
rect 2599 -5618 2641 -5382
rect 2321 -5702 2641 -5618
rect 2321 -5938 2363 -5702
rect 2599 -5938 2641 -5702
rect 2321 -6022 2641 -5938
rect 2321 -6258 2363 -6022
rect 2599 -6258 2641 -6022
rect 2321 -6342 2641 -6258
rect 2321 -6578 2363 -6342
rect 2599 -6578 2641 -6342
rect 2321 -6662 2641 -6578
rect 2321 -6898 2363 -6662
rect 2599 -6898 2641 -6662
rect 2321 -6982 2641 -6898
rect 2321 -7218 2363 -6982
rect 2599 -7218 2641 -6982
rect 2321 -7302 2641 -7218
rect 2321 -7538 2363 -7302
rect 2599 -7538 2641 -7302
rect -239 -7770 81 -7604
rect 2321 -7770 2641 -7538
<< properties >>
string FIXED_BBOX -2619 2640 2461 7720
<< end >>
