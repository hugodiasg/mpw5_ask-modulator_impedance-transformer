magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< metal4 >>
rect -2586 10029 2586 10178
rect -2586 9793 2330 10029
rect 2566 9793 2586 10029
rect -2586 9709 2586 9793
rect -2586 9473 2330 9709
rect 2566 9473 2586 9709
rect -2586 9389 2586 9473
rect -2586 9153 2330 9389
rect 2566 9153 2586 9389
rect -2586 9069 2586 9153
rect -2586 8833 2330 9069
rect 2566 8833 2586 9069
rect -2586 8749 2586 8833
rect -2586 8513 2330 8749
rect 2566 8513 2586 8749
rect -2586 8429 2586 8513
rect -2586 8193 2330 8429
rect 2566 8193 2586 8429
rect -2586 8109 2586 8193
rect -2586 7873 2330 8109
rect 2566 7873 2586 8109
rect -2586 7789 2586 7873
rect -2586 7553 2330 7789
rect 2566 7553 2586 7789
rect -2586 7469 2586 7553
rect -2586 7233 2330 7469
rect 2566 7233 2586 7469
rect -2586 7149 2586 7233
rect -2586 6913 2330 7149
rect 2566 6913 2586 7149
rect -2586 6829 2586 6913
rect -2586 6593 2330 6829
rect 2566 6593 2586 6829
rect -2586 6509 2586 6593
rect -2586 6273 2330 6509
rect 2566 6273 2586 6509
rect -2586 6189 2586 6273
rect -2586 5953 2330 6189
rect 2566 5953 2586 6189
rect -2586 5869 2586 5953
rect -2586 5633 2330 5869
rect 2566 5633 2586 5869
rect -2586 5549 2586 5633
rect -2586 5313 2330 5549
rect 2566 5313 2586 5549
rect -2586 5164 2586 5313
rect -2586 4915 2586 5064
rect -2586 4679 2330 4915
rect 2566 4679 2586 4915
rect -2586 4595 2586 4679
rect -2586 4359 2330 4595
rect 2566 4359 2586 4595
rect -2586 4275 2586 4359
rect -2586 4039 2330 4275
rect 2566 4039 2586 4275
rect -2586 3955 2586 4039
rect -2586 3719 2330 3955
rect 2566 3719 2586 3955
rect -2586 3635 2586 3719
rect -2586 3399 2330 3635
rect 2566 3399 2586 3635
rect -2586 3315 2586 3399
rect -2586 3079 2330 3315
rect 2566 3079 2586 3315
rect -2586 2995 2586 3079
rect -2586 2759 2330 2995
rect 2566 2759 2586 2995
rect -2586 2675 2586 2759
rect -2586 2439 2330 2675
rect 2566 2439 2586 2675
rect -2586 2355 2586 2439
rect -2586 2119 2330 2355
rect 2566 2119 2586 2355
rect -2586 2035 2586 2119
rect -2586 1799 2330 2035
rect 2566 1799 2586 2035
rect -2586 1715 2586 1799
rect -2586 1479 2330 1715
rect 2566 1479 2586 1715
rect -2586 1395 2586 1479
rect -2586 1159 2330 1395
rect 2566 1159 2586 1395
rect -2586 1075 2586 1159
rect -2586 839 2330 1075
rect 2566 839 2586 1075
rect -2586 755 2586 839
rect -2586 519 2330 755
rect 2566 519 2586 755
rect -2586 435 2586 519
rect -2586 199 2330 435
rect 2566 199 2586 435
rect -2586 50 2586 199
rect -2586 -199 2586 -50
rect -2586 -435 2330 -199
rect 2566 -435 2586 -199
rect -2586 -519 2586 -435
rect -2586 -755 2330 -519
rect 2566 -755 2586 -519
rect -2586 -839 2586 -755
rect -2586 -1075 2330 -839
rect 2566 -1075 2586 -839
rect -2586 -1159 2586 -1075
rect -2586 -1395 2330 -1159
rect 2566 -1395 2586 -1159
rect -2586 -1479 2586 -1395
rect -2586 -1715 2330 -1479
rect 2566 -1715 2586 -1479
rect -2586 -1799 2586 -1715
rect -2586 -2035 2330 -1799
rect 2566 -2035 2586 -1799
rect -2586 -2119 2586 -2035
rect -2586 -2355 2330 -2119
rect 2566 -2355 2586 -2119
rect -2586 -2439 2586 -2355
rect -2586 -2675 2330 -2439
rect 2566 -2675 2586 -2439
rect -2586 -2759 2586 -2675
rect -2586 -2995 2330 -2759
rect 2566 -2995 2586 -2759
rect -2586 -3079 2586 -2995
rect -2586 -3315 2330 -3079
rect 2566 -3315 2586 -3079
rect -2586 -3399 2586 -3315
rect -2586 -3635 2330 -3399
rect 2566 -3635 2586 -3399
rect -2586 -3719 2586 -3635
rect -2586 -3955 2330 -3719
rect 2566 -3955 2586 -3719
rect -2586 -4039 2586 -3955
rect -2586 -4275 2330 -4039
rect 2566 -4275 2586 -4039
rect -2586 -4359 2586 -4275
rect -2586 -4595 2330 -4359
rect 2566 -4595 2586 -4359
rect -2586 -4679 2586 -4595
rect -2586 -4915 2330 -4679
rect 2566 -4915 2586 -4679
rect -2586 -5064 2586 -4915
rect -2586 -5313 2586 -5164
rect -2586 -5549 2330 -5313
rect 2566 -5549 2586 -5313
rect -2586 -5633 2586 -5549
rect -2586 -5869 2330 -5633
rect 2566 -5869 2586 -5633
rect -2586 -5953 2586 -5869
rect -2586 -6189 2330 -5953
rect 2566 -6189 2586 -5953
rect -2586 -6273 2586 -6189
rect -2586 -6509 2330 -6273
rect 2566 -6509 2586 -6273
rect -2586 -6593 2586 -6509
rect -2586 -6829 2330 -6593
rect 2566 -6829 2586 -6593
rect -2586 -6913 2586 -6829
rect -2586 -7149 2330 -6913
rect 2566 -7149 2586 -6913
rect -2586 -7233 2586 -7149
rect -2586 -7469 2330 -7233
rect 2566 -7469 2586 -7233
rect -2586 -7553 2586 -7469
rect -2586 -7789 2330 -7553
rect 2566 -7789 2586 -7553
rect -2586 -7873 2586 -7789
rect -2586 -8109 2330 -7873
rect 2566 -8109 2586 -7873
rect -2586 -8193 2586 -8109
rect -2586 -8429 2330 -8193
rect 2566 -8429 2586 -8193
rect -2586 -8513 2586 -8429
rect -2586 -8749 2330 -8513
rect 2566 -8749 2586 -8513
rect -2586 -8833 2586 -8749
rect -2586 -9069 2330 -8833
rect 2566 -9069 2586 -8833
rect -2586 -9153 2586 -9069
rect -2586 -9389 2330 -9153
rect 2566 -9389 2586 -9153
rect -2586 -9473 2586 -9389
rect -2586 -9709 2330 -9473
rect 2566 -9709 2586 -9473
rect -2586 -9793 2586 -9709
rect -2586 -10029 2330 -9793
rect 2566 -10029 2586 -9793
rect -2586 -10178 2586 -10029
<< via4 >>
rect 2330 9793 2566 10029
rect 2330 9473 2566 9709
rect 2330 9153 2566 9389
rect 2330 8833 2566 9069
rect 2330 8513 2566 8749
rect 2330 8193 2566 8429
rect 2330 7873 2566 8109
rect 2330 7553 2566 7789
rect 2330 7233 2566 7469
rect 2330 6913 2566 7149
rect 2330 6593 2566 6829
rect 2330 6273 2566 6509
rect 2330 5953 2566 6189
rect 2330 5633 2566 5869
rect 2330 5313 2566 5549
rect 2330 4679 2566 4915
rect 2330 4359 2566 4595
rect 2330 4039 2566 4275
rect 2330 3719 2566 3955
rect 2330 3399 2566 3635
rect 2330 3079 2566 3315
rect 2330 2759 2566 2995
rect 2330 2439 2566 2675
rect 2330 2119 2566 2355
rect 2330 1799 2566 2035
rect 2330 1479 2566 1715
rect 2330 1159 2566 1395
rect 2330 839 2566 1075
rect 2330 519 2566 755
rect 2330 199 2566 435
rect 2330 -435 2566 -199
rect 2330 -755 2566 -519
rect 2330 -1075 2566 -839
rect 2330 -1395 2566 -1159
rect 2330 -1715 2566 -1479
rect 2330 -2035 2566 -1799
rect 2330 -2355 2566 -2119
rect 2330 -2675 2566 -2439
rect 2330 -2995 2566 -2759
rect 2330 -3315 2566 -3079
rect 2330 -3635 2566 -3399
rect 2330 -3955 2566 -3719
rect 2330 -4275 2566 -4039
rect 2330 -4595 2566 -4359
rect 2330 -4915 2566 -4679
rect 2330 -5549 2566 -5313
rect 2330 -5869 2566 -5633
rect 2330 -6189 2566 -5953
rect 2330 -6509 2566 -6273
rect 2330 -6829 2566 -6593
rect 2330 -7149 2566 -6913
rect 2330 -7469 2566 -7233
rect 2330 -7789 2566 -7553
rect 2330 -8109 2566 -7873
rect 2330 -8429 2566 -8193
rect 2330 -8749 2566 -8513
rect 2330 -9069 2566 -8833
rect 2330 -9389 2566 -9153
rect 2330 -9709 2566 -9473
rect 2330 -10029 2566 -9793
<< mimcap2 >>
rect -2486 10029 2328 10078
rect -2486 5313 -1957 10029
rect 1799 5313 2328 10029
rect -2486 5264 2328 5313
rect -2486 4915 2328 4964
rect -2486 199 -1957 4915
rect 1799 199 2328 4915
rect -2486 150 2328 199
rect -2486 -199 2328 -150
rect -2486 -4915 -1957 -199
rect 1799 -4915 2328 -199
rect -2486 -4964 2328 -4915
rect -2486 -5313 2328 -5264
rect -2486 -10029 -1957 -5313
rect 1799 -10029 2328 -5313
rect -2486 -10078 2328 -10029
<< mimcap2contact >>
rect -1957 5313 1799 10029
rect -1957 199 1799 4915
rect -1957 -4915 1799 -199
rect -1957 -10029 1799 -5313
<< metal5 >>
rect -239 10062 81 10228
rect -1997 10029 1839 10062
rect -1997 5313 -1957 10029
rect 1799 5313 1839 10029
rect -1997 5280 1839 5313
rect 2288 10029 2608 10228
rect 2288 9793 2330 10029
rect 2566 9793 2608 10029
rect 2288 9709 2608 9793
rect 2288 9473 2330 9709
rect 2566 9473 2608 9709
rect 2288 9389 2608 9473
rect 2288 9153 2330 9389
rect 2566 9153 2608 9389
rect 2288 9069 2608 9153
rect 2288 8833 2330 9069
rect 2566 8833 2608 9069
rect 2288 8749 2608 8833
rect 2288 8513 2330 8749
rect 2566 8513 2608 8749
rect 2288 8429 2608 8513
rect 2288 8193 2330 8429
rect 2566 8193 2608 8429
rect 2288 8109 2608 8193
rect 2288 7873 2330 8109
rect 2566 7873 2608 8109
rect 2288 7789 2608 7873
rect 2288 7553 2330 7789
rect 2566 7553 2608 7789
rect 2288 7469 2608 7553
rect 2288 7233 2330 7469
rect 2566 7233 2608 7469
rect 2288 7149 2608 7233
rect 2288 6913 2330 7149
rect 2566 6913 2608 7149
rect 2288 6829 2608 6913
rect 2288 6593 2330 6829
rect 2566 6593 2608 6829
rect 2288 6509 2608 6593
rect 2288 6273 2330 6509
rect 2566 6273 2608 6509
rect 2288 6189 2608 6273
rect 2288 5953 2330 6189
rect 2566 5953 2608 6189
rect 2288 5869 2608 5953
rect 2288 5633 2330 5869
rect 2566 5633 2608 5869
rect 2288 5549 2608 5633
rect 2288 5313 2330 5549
rect 2566 5313 2608 5549
rect -239 4948 81 5280
rect -1997 4915 1839 4948
rect -1997 199 -1957 4915
rect 1799 199 1839 4915
rect -1997 166 1839 199
rect 2288 4915 2608 5313
rect 2288 4679 2330 4915
rect 2566 4679 2608 4915
rect 2288 4595 2608 4679
rect 2288 4359 2330 4595
rect 2566 4359 2608 4595
rect 2288 4275 2608 4359
rect 2288 4039 2330 4275
rect 2566 4039 2608 4275
rect 2288 3955 2608 4039
rect 2288 3719 2330 3955
rect 2566 3719 2608 3955
rect 2288 3635 2608 3719
rect 2288 3399 2330 3635
rect 2566 3399 2608 3635
rect 2288 3315 2608 3399
rect 2288 3079 2330 3315
rect 2566 3079 2608 3315
rect 2288 2995 2608 3079
rect 2288 2759 2330 2995
rect 2566 2759 2608 2995
rect 2288 2675 2608 2759
rect 2288 2439 2330 2675
rect 2566 2439 2608 2675
rect 2288 2355 2608 2439
rect 2288 2119 2330 2355
rect 2566 2119 2608 2355
rect 2288 2035 2608 2119
rect 2288 1799 2330 2035
rect 2566 1799 2608 2035
rect 2288 1715 2608 1799
rect 2288 1479 2330 1715
rect 2566 1479 2608 1715
rect 2288 1395 2608 1479
rect 2288 1159 2330 1395
rect 2566 1159 2608 1395
rect 2288 1075 2608 1159
rect 2288 839 2330 1075
rect 2566 839 2608 1075
rect 2288 755 2608 839
rect 2288 519 2330 755
rect 2566 519 2608 755
rect 2288 435 2608 519
rect 2288 199 2330 435
rect 2566 199 2608 435
rect -239 -166 81 166
rect -1997 -199 1839 -166
rect -1997 -4915 -1957 -199
rect 1799 -4915 1839 -199
rect -1997 -4948 1839 -4915
rect 2288 -199 2608 199
rect 2288 -435 2330 -199
rect 2566 -435 2608 -199
rect 2288 -519 2608 -435
rect 2288 -755 2330 -519
rect 2566 -755 2608 -519
rect 2288 -839 2608 -755
rect 2288 -1075 2330 -839
rect 2566 -1075 2608 -839
rect 2288 -1159 2608 -1075
rect 2288 -1395 2330 -1159
rect 2566 -1395 2608 -1159
rect 2288 -1479 2608 -1395
rect 2288 -1715 2330 -1479
rect 2566 -1715 2608 -1479
rect 2288 -1799 2608 -1715
rect 2288 -2035 2330 -1799
rect 2566 -2035 2608 -1799
rect 2288 -2119 2608 -2035
rect 2288 -2355 2330 -2119
rect 2566 -2355 2608 -2119
rect 2288 -2439 2608 -2355
rect 2288 -2675 2330 -2439
rect 2566 -2675 2608 -2439
rect 2288 -2759 2608 -2675
rect 2288 -2995 2330 -2759
rect 2566 -2995 2608 -2759
rect 2288 -3079 2608 -2995
rect 2288 -3315 2330 -3079
rect 2566 -3315 2608 -3079
rect 2288 -3399 2608 -3315
rect 2288 -3635 2330 -3399
rect 2566 -3635 2608 -3399
rect 2288 -3719 2608 -3635
rect 2288 -3955 2330 -3719
rect 2566 -3955 2608 -3719
rect 2288 -4039 2608 -3955
rect 2288 -4275 2330 -4039
rect 2566 -4275 2608 -4039
rect 2288 -4359 2608 -4275
rect 2288 -4595 2330 -4359
rect 2566 -4595 2608 -4359
rect 2288 -4679 2608 -4595
rect 2288 -4915 2330 -4679
rect 2566 -4915 2608 -4679
rect -239 -5280 81 -4948
rect -1997 -5313 1839 -5280
rect -1997 -10029 -1957 -5313
rect 1799 -10029 1839 -5313
rect -1997 -10062 1839 -10029
rect 2288 -5313 2608 -4915
rect 2288 -5549 2330 -5313
rect 2566 -5549 2608 -5313
rect 2288 -5633 2608 -5549
rect 2288 -5869 2330 -5633
rect 2566 -5869 2608 -5633
rect 2288 -5953 2608 -5869
rect 2288 -6189 2330 -5953
rect 2566 -6189 2608 -5953
rect 2288 -6273 2608 -6189
rect 2288 -6509 2330 -6273
rect 2566 -6509 2608 -6273
rect 2288 -6593 2608 -6509
rect 2288 -6829 2330 -6593
rect 2566 -6829 2608 -6593
rect 2288 -6913 2608 -6829
rect 2288 -7149 2330 -6913
rect 2566 -7149 2608 -6913
rect 2288 -7233 2608 -7149
rect 2288 -7469 2330 -7233
rect 2566 -7469 2608 -7233
rect 2288 -7553 2608 -7469
rect 2288 -7789 2330 -7553
rect 2566 -7789 2608 -7553
rect 2288 -7873 2608 -7789
rect 2288 -8109 2330 -7873
rect 2566 -8109 2608 -7873
rect 2288 -8193 2608 -8109
rect 2288 -8429 2330 -8193
rect 2566 -8429 2608 -8193
rect 2288 -8513 2608 -8429
rect 2288 -8749 2330 -8513
rect 2566 -8749 2608 -8513
rect 2288 -8833 2608 -8749
rect 2288 -9069 2330 -8833
rect 2566 -9069 2608 -8833
rect 2288 -9153 2608 -9069
rect 2288 -9389 2330 -9153
rect 2566 -9389 2608 -9153
rect 2288 -9473 2608 -9389
rect 2288 -9709 2330 -9473
rect 2566 -9709 2608 -9473
rect 2288 -9793 2608 -9709
rect 2288 -10029 2330 -9793
rect 2566 -10029 2608 -9793
rect -239 -10228 81 -10062
rect 2288 -10228 2608 -10029
<< properties >>
string FIXED_BBOX -2586 5164 2428 10178
<< end >>
