magic
tech sky130A
magscale 1 2
timestamp 1647143569
<< pwell >>
rect -268 -1118 268 1118
<< mvnmos >>
rect -50 -870 50 870
<< mvndiff >>
rect -108 833 -50 870
rect -108 799 -96 833
rect -62 799 -50 833
rect -108 765 -50 799
rect -108 731 -96 765
rect -62 731 -50 765
rect -108 697 -50 731
rect -108 663 -96 697
rect -62 663 -50 697
rect -108 629 -50 663
rect -108 595 -96 629
rect -62 595 -50 629
rect -108 561 -50 595
rect -108 527 -96 561
rect -62 527 -50 561
rect -108 493 -50 527
rect -108 459 -96 493
rect -62 459 -50 493
rect -108 425 -50 459
rect -108 391 -96 425
rect -62 391 -50 425
rect -108 357 -50 391
rect -108 323 -96 357
rect -62 323 -50 357
rect -108 289 -50 323
rect -108 255 -96 289
rect -62 255 -50 289
rect -108 221 -50 255
rect -108 187 -96 221
rect -62 187 -50 221
rect -108 153 -50 187
rect -108 119 -96 153
rect -62 119 -50 153
rect -108 85 -50 119
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -119 -50 -85
rect -108 -153 -96 -119
rect -62 -153 -50 -119
rect -108 -187 -50 -153
rect -108 -221 -96 -187
rect -62 -221 -50 -187
rect -108 -255 -50 -221
rect -108 -289 -96 -255
rect -62 -289 -50 -255
rect -108 -323 -50 -289
rect -108 -357 -96 -323
rect -62 -357 -50 -323
rect -108 -391 -50 -357
rect -108 -425 -96 -391
rect -62 -425 -50 -391
rect -108 -459 -50 -425
rect -108 -493 -96 -459
rect -62 -493 -50 -459
rect -108 -527 -50 -493
rect -108 -561 -96 -527
rect -62 -561 -50 -527
rect -108 -595 -50 -561
rect -108 -629 -96 -595
rect -62 -629 -50 -595
rect -108 -663 -50 -629
rect -108 -697 -96 -663
rect -62 -697 -50 -663
rect -108 -731 -50 -697
rect -108 -765 -96 -731
rect -62 -765 -50 -731
rect -108 -799 -50 -765
rect -108 -833 -96 -799
rect -62 -833 -50 -799
rect -108 -870 -50 -833
rect 50 833 108 870
rect 50 799 62 833
rect 96 799 108 833
rect 50 765 108 799
rect 50 731 62 765
rect 96 731 108 765
rect 50 697 108 731
rect 50 663 62 697
rect 96 663 108 697
rect 50 629 108 663
rect 50 595 62 629
rect 96 595 108 629
rect 50 561 108 595
rect 50 527 62 561
rect 96 527 108 561
rect 50 493 108 527
rect 50 459 62 493
rect 96 459 108 493
rect 50 425 108 459
rect 50 391 62 425
rect 96 391 108 425
rect 50 357 108 391
rect 50 323 62 357
rect 96 323 108 357
rect 50 289 108 323
rect 50 255 62 289
rect 96 255 108 289
rect 50 221 108 255
rect 50 187 62 221
rect 96 187 108 221
rect 50 153 108 187
rect 50 119 62 153
rect 96 119 108 153
rect 50 85 108 119
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -119 108 -85
rect 50 -153 62 -119
rect 96 -153 108 -119
rect 50 -187 108 -153
rect 50 -221 62 -187
rect 96 -221 108 -187
rect 50 -255 108 -221
rect 50 -289 62 -255
rect 96 -289 108 -255
rect 50 -323 108 -289
rect 50 -357 62 -323
rect 96 -357 108 -323
rect 50 -391 108 -357
rect 50 -425 62 -391
rect 96 -425 108 -391
rect 50 -459 108 -425
rect 50 -493 62 -459
rect 96 -493 108 -459
rect 50 -527 108 -493
rect 50 -561 62 -527
rect 96 -561 108 -527
rect 50 -595 108 -561
rect 50 -629 62 -595
rect 96 -629 108 -595
rect 50 -663 108 -629
rect 50 -697 62 -663
rect 96 -697 108 -663
rect 50 -731 108 -697
rect 50 -765 62 -731
rect 96 -765 108 -731
rect 50 -799 108 -765
rect 50 -833 62 -799
rect 96 -833 108 -799
rect 50 -870 108 -833
<< mvndiffc >>
rect -96 799 -62 833
rect -96 731 -62 765
rect -96 663 -62 697
rect -96 595 -62 629
rect -96 527 -62 561
rect -96 459 -62 493
rect -96 391 -62 425
rect -96 323 -62 357
rect -96 255 -62 289
rect -96 187 -62 221
rect -96 119 -62 153
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect -96 -153 -62 -119
rect -96 -221 -62 -187
rect -96 -289 -62 -255
rect -96 -357 -62 -323
rect -96 -425 -62 -391
rect -96 -493 -62 -459
rect -96 -561 -62 -527
rect -96 -629 -62 -595
rect -96 -697 -62 -663
rect -96 -765 -62 -731
rect -96 -833 -62 -799
rect 62 799 96 833
rect 62 731 96 765
rect 62 663 96 697
rect 62 595 96 629
rect 62 527 96 561
rect 62 459 96 493
rect 62 391 96 425
rect 62 323 96 357
rect 62 255 96 289
rect 62 187 96 221
rect 62 119 96 153
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
rect 62 -153 96 -119
rect 62 -221 96 -187
rect 62 -289 96 -255
rect 62 -357 96 -323
rect 62 -425 96 -391
rect 62 -493 96 -459
rect 62 -561 96 -527
rect 62 -629 96 -595
rect 62 -697 96 -663
rect 62 -765 96 -731
rect 62 -833 96 -799
<< mvpsubdiff >>
rect -242 1080 242 1092
rect -242 1046 -119 1080
rect -85 1046 -51 1080
rect -17 1046 17 1080
rect 51 1046 85 1080
rect 119 1046 242 1080
rect -242 1034 242 1046
rect -242 969 -184 1034
rect -242 935 -230 969
rect -196 935 -184 969
rect 184 969 242 1034
rect -242 901 -184 935
rect -242 867 -230 901
rect -196 867 -184 901
rect 184 935 196 969
rect 230 935 242 969
rect 184 901 242 935
rect -242 833 -184 867
rect -242 799 -230 833
rect -196 799 -184 833
rect -242 765 -184 799
rect -242 731 -230 765
rect -196 731 -184 765
rect -242 697 -184 731
rect -242 663 -230 697
rect -196 663 -184 697
rect -242 629 -184 663
rect -242 595 -230 629
rect -196 595 -184 629
rect -242 561 -184 595
rect -242 527 -230 561
rect -196 527 -184 561
rect -242 493 -184 527
rect -242 459 -230 493
rect -196 459 -184 493
rect -242 425 -184 459
rect -242 391 -230 425
rect -196 391 -184 425
rect -242 357 -184 391
rect -242 323 -230 357
rect -196 323 -184 357
rect -242 289 -184 323
rect -242 255 -230 289
rect -196 255 -184 289
rect -242 221 -184 255
rect -242 187 -230 221
rect -196 187 -184 221
rect -242 153 -184 187
rect -242 119 -230 153
rect -196 119 -184 153
rect -242 85 -184 119
rect -242 51 -230 85
rect -196 51 -184 85
rect -242 17 -184 51
rect -242 -17 -230 17
rect -196 -17 -184 17
rect -242 -51 -184 -17
rect -242 -85 -230 -51
rect -196 -85 -184 -51
rect -242 -119 -184 -85
rect -242 -153 -230 -119
rect -196 -153 -184 -119
rect -242 -187 -184 -153
rect -242 -221 -230 -187
rect -196 -221 -184 -187
rect -242 -255 -184 -221
rect -242 -289 -230 -255
rect -196 -289 -184 -255
rect -242 -323 -184 -289
rect -242 -357 -230 -323
rect -196 -357 -184 -323
rect -242 -391 -184 -357
rect -242 -425 -230 -391
rect -196 -425 -184 -391
rect -242 -459 -184 -425
rect -242 -493 -230 -459
rect -196 -493 -184 -459
rect -242 -527 -184 -493
rect -242 -561 -230 -527
rect -196 -561 -184 -527
rect -242 -595 -184 -561
rect -242 -629 -230 -595
rect -196 -629 -184 -595
rect -242 -663 -184 -629
rect -242 -697 -230 -663
rect -196 -697 -184 -663
rect -242 -731 -184 -697
rect -242 -765 -230 -731
rect -196 -765 -184 -731
rect -242 -799 -184 -765
rect -242 -833 -230 -799
rect -196 -833 -184 -799
rect -242 -867 -184 -833
rect -242 -901 -230 -867
rect -196 -901 -184 -867
rect 184 867 196 901
rect 230 867 242 901
rect 184 833 242 867
rect 184 799 196 833
rect 230 799 242 833
rect 184 765 242 799
rect 184 731 196 765
rect 230 731 242 765
rect 184 697 242 731
rect 184 663 196 697
rect 230 663 242 697
rect 184 629 242 663
rect 184 595 196 629
rect 230 595 242 629
rect 184 561 242 595
rect 184 527 196 561
rect 230 527 242 561
rect 184 493 242 527
rect 184 459 196 493
rect 230 459 242 493
rect 184 425 242 459
rect 184 391 196 425
rect 230 391 242 425
rect 184 357 242 391
rect 184 323 196 357
rect 230 323 242 357
rect 184 289 242 323
rect 184 255 196 289
rect 230 255 242 289
rect 184 221 242 255
rect 184 187 196 221
rect 230 187 242 221
rect 184 153 242 187
rect 184 119 196 153
rect 230 119 242 153
rect 184 85 242 119
rect 184 51 196 85
rect 230 51 242 85
rect 184 17 242 51
rect 184 -17 196 17
rect 230 -17 242 17
rect 184 -51 242 -17
rect 184 -85 196 -51
rect 230 -85 242 -51
rect 184 -119 242 -85
rect 184 -153 196 -119
rect 230 -153 242 -119
rect 184 -187 242 -153
rect 184 -221 196 -187
rect 230 -221 242 -187
rect 184 -255 242 -221
rect 184 -289 196 -255
rect 230 -289 242 -255
rect 184 -323 242 -289
rect 184 -357 196 -323
rect 230 -357 242 -323
rect 184 -391 242 -357
rect 184 -425 196 -391
rect 230 -425 242 -391
rect 184 -459 242 -425
rect 184 -493 196 -459
rect 230 -493 242 -459
rect 184 -527 242 -493
rect 184 -561 196 -527
rect 230 -561 242 -527
rect 184 -595 242 -561
rect 184 -629 196 -595
rect 230 -629 242 -595
rect 184 -663 242 -629
rect 184 -697 196 -663
rect 230 -697 242 -663
rect 184 -731 242 -697
rect 184 -765 196 -731
rect 230 -765 242 -731
rect 184 -799 242 -765
rect 184 -833 196 -799
rect 230 -833 242 -799
rect 184 -867 242 -833
rect -242 -935 -184 -901
rect -242 -969 -230 -935
rect -196 -969 -184 -935
rect 184 -901 196 -867
rect 230 -901 242 -867
rect 184 -935 242 -901
rect -242 -1034 -184 -969
rect 184 -969 196 -935
rect 230 -969 242 -935
rect 184 -1034 242 -969
rect -242 -1046 242 -1034
rect -242 -1080 -119 -1046
rect -85 -1080 -51 -1046
rect -17 -1080 17 -1046
rect 51 -1080 85 -1046
rect 119 -1080 242 -1046
rect -242 -1092 242 -1080
<< mvpsubdiffcont >>
rect -119 1046 -85 1080
rect -51 1046 -17 1080
rect 17 1046 51 1080
rect 85 1046 119 1080
rect -230 935 -196 969
rect -230 867 -196 901
rect 196 935 230 969
rect -230 799 -196 833
rect -230 731 -196 765
rect -230 663 -196 697
rect -230 595 -196 629
rect -230 527 -196 561
rect -230 459 -196 493
rect -230 391 -196 425
rect -230 323 -196 357
rect -230 255 -196 289
rect -230 187 -196 221
rect -230 119 -196 153
rect -230 51 -196 85
rect -230 -17 -196 17
rect -230 -85 -196 -51
rect -230 -153 -196 -119
rect -230 -221 -196 -187
rect -230 -289 -196 -255
rect -230 -357 -196 -323
rect -230 -425 -196 -391
rect -230 -493 -196 -459
rect -230 -561 -196 -527
rect -230 -629 -196 -595
rect -230 -697 -196 -663
rect -230 -765 -196 -731
rect -230 -833 -196 -799
rect -230 -901 -196 -867
rect 196 867 230 901
rect 196 799 230 833
rect 196 731 230 765
rect 196 663 230 697
rect 196 595 230 629
rect 196 527 230 561
rect 196 459 230 493
rect 196 391 230 425
rect 196 323 230 357
rect 196 255 230 289
rect 196 187 230 221
rect 196 119 230 153
rect 196 51 230 85
rect 196 -17 230 17
rect 196 -85 230 -51
rect 196 -153 230 -119
rect 196 -221 230 -187
rect 196 -289 230 -255
rect 196 -357 230 -323
rect 196 -425 230 -391
rect 196 -493 230 -459
rect 196 -561 230 -527
rect 196 -629 230 -595
rect 196 -697 230 -663
rect 196 -765 230 -731
rect 196 -833 230 -799
rect -230 -969 -196 -935
rect 196 -901 230 -867
rect 196 -969 230 -935
rect -119 -1080 -85 -1046
rect -51 -1080 -17 -1046
rect 17 -1080 51 -1046
rect 85 -1080 119 -1046
<< poly >>
rect -50 942 50 958
rect -50 908 -17 942
rect 17 908 50 942
rect -50 870 50 908
rect -50 -908 50 -870
rect -50 -942 -17 -908
rect 17 -942 50 -908
rect -50 -958 50 -942
<< polycont >>
rect -17 908 17 942
rect -17 -942 17 -908
<< locali >>
rect -230 1046 -161 1080
rect -127 1046 -119 1080
rect -55 1046 -51 1080
rect 51 1046 55 1080
rect 119 1046 127 1080
rect 161 1046 230 1080
rect -230 969 -196 1046
rect 196 969 230 1046
rect -230 901 -196 935
rect -50 908 -17 942
rect 17 908 50 942
rect 196 901 230 935
rect -230 833 -196 867
rect -230 765 -196 799
rect -230 697 -196 731
rect -230 629 -196 663
rect -230 561 -196 595
rect -230 493 -196 527
rect -230 425 -196 459
rect -230 357 -196 391
rect -230 289 -196 323
rect -230 221 -196 255
rect -230 153 -196 187
rect -230 85 -196 119
rect -230 17 -196 51
rect -230 -51 -196 -17
rect -230 -119 -196 -85
rect -230 -187 -196 -153
rect -230 -255 -196 -221
rect -230 -323 -196 -289
rect -230 -391 -196 -357
rect -230 -459 -196 -425
rect -230 -527 -196 -493
rect -230 -595 -196 -561
rect -230 -663 -196 -629
rect -230 -731 -196 -697
rect -230 -799 -196 -765
rect -230 -867 -196 -833
rect -96 833 -62 874
rect -96 765 -62 799
rect -96 697 -62 731
rect -96 629 -62 631
rect -96 593 -62 595
rect -96 521 -62 527
rect -96 449 -62 459
rect -96 377 -62 391
rect -96 305 -62 323
rect -96 233 -62 255
rect -96 161 -62 187
rect -96 89 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -89
rect -96 -187 -62 -161
rect -96 -255 -62 -233
rect -96 -323 -62 -305
rect -96 -391 -62 -377
rect -96 -459 -62 -449
rect -96 -527 -62 -521
rect -96 -595 -62 -593
rect -96 -631 -62 -629
rect -96 -731 -62 -697
rect -96 -799 -62 -765
rect -96 -874 -62 -833
rect 62 833 96 874
rect 62 765 96 799
rect 62 697 96 731
rect 62 629 96 631
rect 62 593 96 595
rect 62 521 96 527
rect 62 449 96 459
rect 62 377 96 391
rect 62 305 96 323
rect 62 233 96 255
rect 62 161 96 187
rect 62 89 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -89
rect 62 -187 96 -161
rect 62 -255 96 -233
rect 62 -323 96 -305
rect 62 -391 96 -377
rect 62 -459 96 -449
rect 62 -527 96 -521
rect 62 -595 96 -593
rect 62 -631 96 -629
rect 62 -731 96 -697
rect 62 -799 96 -765
rect 62 -874 96 -833
rect 196 833 230 867
rect 196 765 230 799
rect 196 697 230 731
rect 196 629 230 663
rect 196 561 230 595
rect 196 493 230 527
rect 196 425 230 459
rect 196 357 230 391
rect 196 289 230 323
rect 196 221 230 255
rect 196 153 230 187
rect 196 85 230 119
rect 196 17 230 51
rect 196 -51 230 -17
rect 196 -119 230 -85
rect 196 -187 230 -153
rect 196 -255 230 -221
rect 196 -323 230 -289
rect 196 -391 230 -357
rect 196 -459 230 -425
rect 196 -527 230 -493
rect 196 -595 230 -561
rect 196 -663 230 -629
rect 196 -731 230 -697
rect 196 -799 230 -765
rect 196 -867 230 -833
rect -230 -935 -196 -901
rect -50 -942 -17 -908
rect 17 -942 50 -908
rect 196 -935 230 -901
rect -230 -1046 -196 -969
rect 196 -1046 230 -969
rect -230 -1080 -119 -1046
rect -85 -1080 -51 -1046
rect -17 -1080 17 -1046
rect 51 -1080 85 -1046
rect 119 -1080 230 -1046
<< viali >>
rect -161 1046 -127 1080
rect -89 1046 -85 1080
rect -85 1046 -55 1080
rect -17 1046 17 1080
rect 55 1046 85 1080
rect 85 1046 89 1080
rect 127 1046 161 1080
rect -17 908 17 942
rect -96 663 -62 665
rect -96 631 -62 663
rect -96 561 -62 593
rect -96 559 -62 561
rect -96 493 -62 521
rect -96 487 -62 493
rect -96 425 -62 449
rect -96 415 -62 425
rect -96 357 -62 377
rect -96 343 -62 357
rect -96 289 -62 305
rect -96 271 -62 289
rect -96 221 -62 233
rect -96 199 -62 221
rect -96 153 -62 161
rect -96 127 -62 153
rect -96 85 -62 89
rect -96 55 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -55
rect -96 -89 -62 -85
rect -96 -153 -62 -127
rect -96 -161 -62 -153
rect -96 -221 -62 -199
rect -96 -233 -62 -221
rect -96 -289 -62 -271
rect -96 -305 -62 -289
rect -96 -357 -62 -343
rect -96 -377 -62 -357
rect -96 -425 -62 -415
rect -96 -449 -62 -425
rect -96 -493 -62 -487
rect -96 -521 -62 -493
rect -96 -561 -62 -559
rect -96 -593 -62 -561
rect -96 -663 -62 -631
rect -96 -665 -62 -663
rect 62 663 96 665
rect 62 631 96 663
rect 62 561 96 593
rect 62 559 96 561
rect 62 493 96 521
rect 62 487 96 493
rect 62 425 96 449
rect 62 415 96 425
rect 62 357 96 377
rect 62 343 96 357
rect 62 289 96 305
rect 62 271 96 289
rect 62 221 96 233
rect 62 199 96 221
rect 62 153 96 161
rect 62 127 96 153
rect 62 85 96 89
rect 62 55 96 85
rect 62 -17 96 17
rect 62 -85 96 -55
rect 62 -89 96 -85
rect 62 -153 96 -127
rect 62 -161 96 -153
rect 62 -221 96 -199
rect 62 -233 96 -221
rect 62 -289 96 -271
rect 62 -305 96 -289
rect 62 -357 96 -343
rect 62 -377 96 -357
rect 62 -425 96 -415
rect 62 -449 96 -425
rect 62 -493 96 -487
rect 62 -521 96 -493
rect 62 -561 96 -559
rect 62 -593 96 -561
rect 62 -663 96 -631
rect 62 -665 96 -663
rect -17 -942 17 -908
<< metal1 >>
rect -208 1080 208 1086
rect -208 1046 -161 1080
rect -127 1046 -89 1080
rect -55 1046 -17 1080
rect 17 1046 55 1080
rect 89 1046 127 1080
rect 161 1046 208 1080
rect -208 1040 208 1046
rect -46 942 46 948
rect -46 908 -17 942
rect 17 908 46 942
rect -46 902 46 908
rect -102 665 -56 698
rect -102 631 -96 665
rect -62 631 -56 665
rect -102 593 -56 631
rect -102 559 -96 593
rect -62 559 -56 593
rect -102 521 -56 559
rect -102 487 -96 521
rect -62 487 -56 521
rect -102 449 -56 487
rect -102 415 -96 449
rect -62 415 -56 449
rect -102 377 -56 415
rect -102 343 -96 377
rect -62 343 -56 377
rect -102 305 -56 343
rect -102 271 -96 305
rect -62 271 -56 305
rect -102 233 -56 271
rect -102 199 -96 233
rect -62 199 -56 233
rect -102 161 -56 199
rect -102 127 -96 161
rect -62 127 -56 161
rect -102 89 -56 127
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -127 -56 -89
rect -102 -161 -96 -127
rect -62 -161 -56 -127
rect -102 -199 -56 -161
rect -102 -233 -96 -199
rect -62 -233 -56 -199
rect -102 -271 -56 -233
rect -102 -305 -96 -271
rect -62 -305 -56 -271
rect -102 -343 -56 -305
rect -102 -377 -96 -343
rect -62 -377 -56 -343
rect -102 -415 -56 -377
rect -102 -449 -96 -415
rect -62 -449 -56 -415
rect -102 -487 -56 -449
rect -102 -521 -96 -487
rect -62 -521 -56 -487
rect -102 -559 -56 -521
rect -102 -593 -96 -559
rect -62 -593 -56 -559
rect -102 -631 -56 -593
rect -102 -665 -96 -631
rect -62 -665 -56 -631
rect -102 -698 -56 -665
rect 56 665 102 698
rect 56 631 62 665
rect 96 631 102 665
rect 56 593 102 631
rect 56 559 62 593
rect 96 559 102 593
rect 56 521 102 559
rect 56 487 62 521
rect 96 487 102 521
rect 56 449 102 487
rect 56 415 62 449
rect 96 415 102 449
rect 56 377 102 415
rect 56 343 62 377
rect 96 343 102 377
rect 56 305 102 343
rect 56 271 62 305
rect 96 271 102 305
rect 56 233 102 271
rect 56 199 62 233
rect 96 199 102 233
rect 56 161 102 199
rect 56 127 62 161
rect 96 127 102 161
rect 56 89 102 127
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -127 102 -89
rect 56 -161 62 -127
rect 96 -161 102 -127
rect 56 -199 102 -161
rect 56 -233 62 -199
rect 96 -233 102 -199
rect 56 -271 102 -233
rect 56 -305 62 -271
rect 96 -305 102 -271
rect 56 -343 102 -305
rect 56 -377 62 -343
rect 96 -377 102 -343
rect 56 -415 102 -377
rect 56 -449 62 -415
rect 96 -449 102 -415
rect 56 -487 102 -449
rect 56 -521 62 -487
rect 96 -521 102 -487
rect 56 -559 102 -521
rect 56 -593 62 -559
rect 96 -593 102 -559
rect 56 -631 102 -593
rect 56 -665 62 -631
rect 96 -665 102 -631
rect 56 -698 102 -665
rect -46 -908 46 -902
rect -46 -942 -17 -908
rect 17 -942 46 -908
rect -46 -948 46 -942
<< properties >>
string FIXED_BBOX -212 -1062 212 1062
<< end >>
